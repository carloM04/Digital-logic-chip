-- TB EXAMPLE PFRL 2024-2025

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity tb_gen2_mod5 is
end tb_gen2_mod5;

architecture project_tb_arch of tb_gen2_mod5 is

    constant CLOCK_PERIOD : time := 20 ns;

    -- Signals to be connected to the component
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);

    -- Signals for the memory
    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    -- Memory
    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

    -- Scenario
    type scenario_config_type is array (0 to 16) of integer;
    constant SCENARIO_LENGTH : integer := 2000;
    constant SCENARIO_LENGTH_STL : std_logic_vector(15 downto 0) := std_logic_vector(to_unsigned(SCENARIO_LENGTH, 16));
    type scenario_type is array (0 to SCENARIO_LENGTH-1) of integer;

    signal scenario_config : scenario_config_type := (to_integer(unsigned(SCENARIO_LENGTH_STL(15 downto 8))),   -- K1
                                                      to_integer(unsigned(SCENARIO_LENGTH_STL(7 downto 0))),    -- K2
                                                      1,                                                        -- S
                                                      11, -3, 5, 9, -4, 5, 10, -9, -10, -1, 21, -1, 3, 5           -- C1-C14
                                                      );
    signal scenario_input : scenario_type := (69, -113, -79, -87, 92, -68, 57, 71, 39, -10, -37, -23, -100, 0, 21, -100, 10, -112, 15, 82, 33, -105, 62, -56, -123, 8, -121, 39, -69, 72, 89, 52, 126, -60, -105, 121, 35, -100, -18, 72, -91, -43, -111, 46, -123, 12, -35, -55, 99, -47, -128, 85, 9, -6, 83, -39, -30, 0, -35, -63, 37, 111, 11, 103, -24, -60, -63, 57, -74, 98, -12, -76, 88, 52, -123, 23, 61, 102, 44, 56, 99, 90, 3, 105, 82, 106, 83, 6, -1, -39, -45, -26, 69, 51, 77, -54, 94, 82, 34, -47, -7, 82, -78, -5, 18, -73, -106, -41, 97, -32, -71, -96, 99, -7, -109, -123, -78, -76, 36, -105, 122, 117, 19, -18, 121, 35, -6, 100, -52, 111, 30, 17, -55, -7, -44, -18, -32, -10, 35, -40, -77, 92, -77, 58, 42, -31, 19, 52, -12, -36, -41, -93, -59, -123, 1, 122, -108, 30, 22, -55, -3, 9, 3, -95, -120, 69, 54, 103, -8, -80, 3, 85, -33, -39, 77, 119, -50, 101, 61, -68, -70, -84, 42, 109, -30, -59, 5, 15, -4, -93, 19, -33, 83, -122, 72, -69, 69, 10, 82, 33, 51, -17, 106, -95, -86, -63, -14, -46, -100, -113, -100, 58, -76, -25, 59, -14, 20, 38, -62, -110, 62, 123, -11, 43, 78, -26, 79, 91, 23, -58, -46, 64, 100, 64, 107, -52, -90, 117, 86, 80, -61, -88, -62, 39, -38, -40, -39, -21, -80, -44, 2, 100, -14, -63, -124, 9, -121, -68, -19, 11, -75, 10, -27, 123, 114, -37, -7, 79, 98, 119, -29, -22, -97, -75, 67, 42, -9, -127, -83, -13, -34, 57, -57, 58, -23, -121, 50, 70, 102, 5, 102, -55, 99, 17, 47, -123, 77, 119, 59, 32, 99, -4, -39, -42, -92, 53, -95, 48, 33, -120, 94, 32, 36, 48, 72, -50, -107, -67, 126, 29, -26, 27, 62, 57, -13, -48, 33, 21, 102, 36, 22, -92, 10, -18, -9, 98, 0, 25, -73, -31, -3, 62, 29, -105, -25, 51, -99, -48, -44, 116, -111, 84, 83, 46, -64, 111, 26, -101, -1, 60, 89, 72, 125, -40, 56, -92, 114, 21, 29, -98, -17, -31, -127, -99, -80, -24, 13, -100, -88, 50, 37, 53, 61, -94, -15, -55, -15, -74, 87, -12, -75, 78, 2, 98, -60, -105, 34, 120, 104, 57, 19, 21, -69, 46, 10, -66, 91, 43, 64, 54, -35, -92, 60, -36, -41, 27, 75, 93, 15, 42, 68, 109, 122, -126, 38, -54, 82, -13, 100, 50, -12, 72, 127, -103, 48, -41, 124, 20, 46, 49, 68, -30, -121, -37, 89, 105, -38, -61, -88, -51, -52, -125, -113, -40, -34, -116, 63, 124, 59, -21, 120, 121, 47, 65, 88, 15, 78, -60, -29, 92, -60, -36, -98, -51, -66, 48, -68, 86, 95, 122, 10, -68, -21, -23, 97, -111, 67, -23, -50, -65, -15, -44, 26, -70, 24, 49, -73, -124, -116, -14, 5, -113, -13, -109, -80, 48, -29, 47, -94, -50, -52, 25, -88, -89, 38, 30, -97, -116, 20, 42, 11, -66, -56, -96, -102, -11, 114, 20, -57, -20, 81, 10, 63, -30, -94, -56, -36, -17, 105, -111, 127, -103, -29, -60, 102, 51, 0, -105, -59, 20, 78, 0, -69, 75, 0, 123, 50, 113, 92, -36, -125, -123, -20, -61, -105, -102, 28, -40, -119, -14, -45, -118, 105, 45, 20, -9, -40, 12, 100, 9, -26, 3, 84, -22, -30, 64, 42, -41, 28, -90, 38, -65, 99, -10, -23, 21, -1, -102, -68, 30, -30, 42, -21, -92, 40, -98, 22, -29, 110, -67, 55, -53, 111, 12, 19, -21, -10, 120, 17, 78, 8, 7, -81, 25, 73, 67, 50, 57, 16, -85, -113, -85, -40, -24, 32, -114, -21, 71, -29, -37, 59, 103, -96, 15, 101, -20, -77, 80, 52, -44, -78, 125, -21, 70, -38, -24, -83, 78, 30, 32, -65, -90, 28, -128, -18, -38, -71, 63, -103, 12, 112, -109, -34, 115, -24, 66, -73, -101, 69, -53, 14, -53, -124, -48, 122, -110, 94, 45, -20, -63, 52, -3, -30, -97, 73, 57, 110, -45, 97, 76, 23, 70, 19, -118, 19, -82, 52, 68, 57, -53, 58, -91, -91, -19, -98, -24, 24, 110, 80, -82, -23, 44, -118, -29, -22, 49, 61, -121, -18, -85, 105, 107, 73, 44, 60, -126, 32, 29, -27, 68, 10, -128, 0, 96, -2, -4, -32, -108, 71, 2, 21, 86, 41, 74, -46, -115, 3, 0, -105, -21, -21, 84, -7, -29, -88, -82, 29, -34, -28, -10, -123, -1, -110, -2, -97, -65, -47, -41, -85, -3, -99, 24, -124, -71, 38, -96, 75, 30, -97, -16, 54, -54, 99, -25, 33, 100, -112, -3, -55, -2, -25, 125, 63, 28, 59, 96, 122, -86, -115, 22, -10, -23, -119, 98, 97, 9, -68, 92, 34, 34, -37, 79, -24, 125, 18, 28, -14, 19, -76, -49, -90, 37, 64, -33, -123, 64, 69, -63, 51, -103, -79, 97, 53, -95, 107, -45, 73, 97, 82, 108, -69, 108, -60, -102, 101, 52, -79, 14, -12, -4, 123, -59, -1, -79, -30, 31, 102, 106, -54, -16, -28, 77, 90, 108, 72, 91, 30, -9, -50, 113, -17, -49, 28, 23, -108, -109, 106, -113, -22, 41, -77, -33, -27, 9, -127, -27, 10, -5, 102, 120, -67, -88, 29, -114, -37, -16, -32, 90, 88, 4, 93, -102, -107, -15, -6, 33, -107, -117, 64, -59, -128, -85, -123, -88, -19, 41, 123, 87, -122, -54, -109, 70, -79, -96, 31, -115, -100, 61, -118, 48, 112, 118, -105, 80, 52, -97, -92, -120, -97, 56, 112, 29, -114, -50, 111, 109, -59, 75, 50, -5, -34, -7, -11, -39, 84, -106, 10, 24, 97, -99, 42, -49, 51, 7, -23, 75, -113, 52, -81, -102, 57, 105, 86, 63, 74, -9, -113, -89, -52, 9, 108, -2, 39, 87, 15, 27, -13, -13, 5, 25, 108, 67, -90, -2, -125, -87, 95, -69, -13, 125, 89, 100, 29, 71, -61, 114, -3, 6, 82, -105, -18, 54, -22, 119, 22, 60, 14, 84, 18, -79, 124, -120, 119, 89, 4, -24, 127, -8, -72, -54, -116, 77, -20, 45, 61, 115, 60, 55, 104, 124, 82, -4, -97, -103, -9, -7, 14, 125, -118, 70, 38, -109, -37, 22, -54, 122, 38, -90, -8, 46, -93, -12, 8, 11, 51, 48, 10, 60, -66, -61, -101, -126, 51, -18, 23, 73, 116, -94, -95, 121, -58, 107, 71, -115, -122, 126, 100, 104, 82, 81, 56, -93, 112, -41, -34, -96, -77, 30, -114, -28, 63, 72, -21, 59, -42, 80, 39, 14, -103, -102, 88, -99, -16, 55, -18, -108, 107, -116, -100, -104, 59, -111, -101, 122, 50, 83, 36, -48, 54, 53, -58, 23, -85, 37, -58, -69, -68, -87, -47, -116, -49, -108, 123, 8, 2, 120, 94, -97, 26, 105, 17, 71, 95, 125, -111, -111, 54, 114, 116, -100, 56, -51, -108, 72, -25, 88, 95, 126, 60, -77, -108, 72, 20, -84, -55, -128, 17, -6, 67, 1, 127, 5, 120, 30, -128, -96, -38, 12, 99, 65, -22, -8, -114, 35, -91, 16, 126, -57, -26, -44, 65, -3, -52, -32, -110, -48, -34, -42, -68, 71, -113, -119, 109, -102, -6, -31, 27, -45, 47, 100, 44, 31, -75, 95, 20, 42, -128, -116, -80, 115, 105, -28, -51, -84, 19, 127, -76, 12, -104, 34, -20, -1, -109, -127, 76, 17, -4, 58, 116, -24, -69, 71, -54, -37, -65, 23, -19, 101, 12, -60, -86, -15, -121, 13, 85, 117, -60, -42, 16, -13, -21, -36, -61, -38, -109, 32, -45, 25, -119, 18, 75, 101, -68, -120, -92, 36, -41, -23, 80, -45, -29, -126, -124, 109, 61, -62, -7, -16, 48, 30, -12, 123, 10, 23, 76, -24, 15, -50, -44, -125, 30, -114, -92, 110, -8, -23, 79, 69, -35, 52, -32, 87, -98, -58, 39, 117, -111, 105, -103, -85, 100, 0, -125, 13, 34, -15, 13, -114, -111, 123, -97, -91, 86, -25, -28, -43, 87, -52, -114, 115, 2, 85, -103, -127, 113, 105, 105, 31, 7, -124, -37, 34, -82, -80, -23, -86, 67, -41, -114, -127, -32, -52, 43, -72, -11, -86, 104, 42, 77, -124, 60, 124, -125, 41, -75, 80, 16, 113, -87, 110, 123, 15, 58, -30, -52, 108, -106, 110, -14, 83, 64, -66, -39, 11, 107, -95, 60, 73, -40, -128, 127, -74, 83, -79, 79, 56, 68, -96, 43, -104, 100, 124, -52, -25, 44, 52, 2, 20, -53, -55, -4, 19, 103, -50, 94, -42, 94, 99, 107, -108, 18, -68, 28, 106, -58, -86, -15, 3, 91, 7, -79, -125, 86, 62, 91, 89, 73, 2, -117, -55, 12, -107, -117, 15, -36, 9, 71, 29, 100, 94, -6, -46, 85, 51, -28, 119, -118, 65, -81, 57, -103, 100, 71, 74, 93, -108, -98, -49, 71, -128, 77, 9, -90, 44, 26, -29, -40, -47, -2, -27, 33, -65, -30, -57, -85, 70, 47, -101, 25, 49, 118, -52, 77, -13, -91, 45, 43, -127, -95, -45, -111, 83, -66, -38, -74, 13, 35, -94, -35, -64, -17, -121, -90, 4, 44, 105, 35, 56, -118, -64, 52, -126, 14, -73, 69, 45, 115, 17, -28, 4, -72, -99, 43, -80, 121, 94, 92, -6, -55, 26, 85, 81, -109, 22, -121, 79, 8, 42, 76, 83, 8, -116, -14, 78, 70, -64, -49, 101, 114, 36, 21, -43, -38, 81, 78, -56, -87, 59, 34, 39, -115, 5, -119, -65, -102, -84, -89, 24, -83, -111, 15, 119, -80, -74, -60, -92, -87, -82, 74, 52, -118, 41, -7, -75, 44, 121, -95, -33, 34, 32, 89, 11, -92, 123, -110, 84, 56, -49, 63, 22, 52, -39, 127, 64, -49, -128, -92, -58, 103, -92, 101, 55, -46, -92, 99, 88, -2, -42, -70, -35, 74, -1, 43, -93, -111, 103, -104, -113, 6, 1, 61, -1, -88, 62, -21, -20, 1, 4, 76, 63, -26, -15, 69, 21, -75, 53, 111, -70, -96, 99, -101, -83, -10, -20, -56, -18, 121, -82, -31, 9, -125, 112, -117, 49, 58, -72, 11, 4, 111, 107, -107, 119, -28, -34, -47, -36, 105, 21, 73, 48, 92, 34, -17, -125, 62, -40, -100, 11, -104, 57, -87, 64, 111, 28, 28, -61, -69, 96, -6, 85, -69, 107, -27, 38, 34, -24, 59, 56, -45, 100, -34, -66, 127, -60, -127, -72, -13, -106, -41, -41, 111, 66, -23, -87, -80, -12, 90, 86, 110, -94, -34, 46, -87, -85, -41, 72, 59, 66, -6, -20, 82, 69, 108, -7, -46, -72, 8, 124, -14, 93, -77, 77, 49, -89, 40, -12, -11, -40, -108, -82, -19, -104, 13, 121, 51, 80, 125, -7, -46, 100, 73, -80, 63, 74, 37, 67, -52, 81, 13, -93, -35, 63, 74, 77, 35, 76, 33, -66, 18, 11, 39, -111, -122, 27, 11, 71, 36, -77, 76, -102, 74, 93, -77, 76, 41, -23, 38, -44, -70, -40, -63, -126, 117, -81, 98, -51, 102, -25, -46, -18, -60, -40, -46, -3, 24, -67, 23, 56, -9, -80, 61, 22, -17, 86, 18, -20, -16, -49, -13, 46, -92, -124, -48, 127, -61, -34, -80, 29, 102, 28, -92, -72, 106, 39, 41, -29, 70, 118, -76, -46, -69, -3, 6, 115, -20, -103, 64, -89, 36, 33, 85, 81, 85, -17, 61, -41, -13, -23, 74, 127, 25, 75, 18, -5, 35, -4, -100, -20, 28, 88, 97, 91, 43, 127, 123, -83, 100, 110, -66, -46, 23, -93, 5, 50, 18, 123, -13, 96, -73, 45, 95, 87, 29, -59, -56, 66, -26, -74, -14, 64, 7, 19, 17, 74, 83, -29, -120, -119, -58, 114, -25, 64, 82, 80, -6, -127, 75, -32, -6, -55, -98, -12, 70, -109, -50, -114, 18, -124, 58, -68, -92, -77, -84, -4, 86, 49, -12, -17, -62, -83);

    signal scenario_output : scenario_type :=(13, -35, -36, -20, 73, 6, 18, 17, 8, -32, -34, -7, -34, 6, 20, -24, 10, -19, 11, 44, 24, -66, 1, -14, -39, 2, -10, 44, 1, 48, 35, 1, 22, -34, -72, 27, 42, -42, -37, 26, -15, -28, -39, 38, -24, 20, 2, -15, 40, 3, -53, 30, 30, -2, 13, -17, -28, -4, 10, -10, 26, 56, -2, 3, -25, -41, -28, 39, -14, 38, 7, -40, 13, 39, -35, -3, 38, 58, 10, -3, 18, 25, -13, 17, 14, 15, -5, -34, -32, -21, -7, 5, 36, 30, 30, -32, 9, 20, 9, -46, -24, 32, -24, -25, 0, -5, -35, -11, 51, 13, -27, -52, 36, 10, -47, -54, -10, 14, 61, -7, 46, 59, 8, -44, 28, 10, -14, 19, -22, 19, -1, -7, -43, -10, -10, 6, -3, -2, 24, -8, -30, 41, -10, 17, 18, -7, -12, 11, -11, -31, -30, -28, 5, -22, 20, 76, -24, -10, 7, -7, -15, -5, 10, -23, -31, 44, 42, 37, -14, -51, -17, 48, 12, -26, 23, 61, -29, -5, 0, -32, -35, -23, 28, 59, -3, -43, -15, 15, 5, -29, 1, 2, 39, -39, 23, -10, 37, 7, 27, 4, 0, -37, 14, -42, -46, -30, 10, -4, -20, -29, -15, 59, 7, -2, 28, 5, -11, 6, -7, -41, 28, 77, 1, -9, 21, -10, 3, 15, 1, -35, -22, 39, 49, 4, 15, -30, -47, 31, 38, 11, -52, -55, -27, 32, 6, -17, -19, 4, -5, 0, 9, 40, -4, -45, -65, 13, -10, -9, 9, 32, -4, 21, 1, 47, 46, -18, -25, 18, 34, 19, -49, -37, -38, -15, 31, 26, -6, -62, -27, 17, 21, 36, -24, 14, 2, -30, 18, 53, 43, -14, 14, -32, 9, -2, 23, -51, 21, 61, 27, -25, 0, -25, -34, -30, -25, 39, -21, 24, 27, -32, 26, 31, 12, -14, 3, -22, -45, -26, 70, 41, -12, -12, 14, 18, -14, -25, 12, 18, 29, -1, -11, -55, 3, 9, 9, 30, -3, -6, -34, -7, 0, 29, 18, -52, -29, 26, -6, -22, -5, 76, -19, 13, 32, 25, -57, 13, 17, -34, -9, 45, 46, 13, 13, -37, -2, -42, 30, 5, 2, -66, -25, -7, -29, -23, -7, 14, 34, -11, -21, 40, 35, 14, 2, -51, -27, -8, 15, -22, 44, 13, -22, 17, 0, 30, -20, -37, 15, 70, 45, -11, -28, -12, -41, 14, 20, -13, 30, 21, 5, -1, -27, -55, 20, 14, 1, 11, 40, 39, 0, 2, 0, 22, 22, -70, -17, -9, 51, -2, 34, 19, -22, -1, 38, -40, -4, -13, 56, 11, 1, -18, 3, -18, -45, -14, 46, 48, -30, -56, -51, -14, 0, -23, -30, 15, 41, -5, 34, 74, 41, -29, 19, 44, 2, -9, 2, -20, 9, -37, -30, 21, -17, -28, -35, -3, 2, 54, 7, 38, 27, 30, -28, -51, -29, 0, 51, -39, 4, -8, -14, -27, 3, 1, 27, -19, -2, 9, -24, -52, -41, 21, 31, -30, 0, -18, -5, 32, 8, 14, -35, -24, -20, 31, -8, -32, 10, 35, -20, -46, 14, 39, 7, -44, -30, -11, -6, 15, 65, 28, -31, -21, 35, 3, 2, -28, -45, -13, 4, 21, 49, -41, 25, -28, -2, -21, 46, 20, -7, -51, -22, 18, 54, 8, -30, 25, 19, 53, 3, 4, -11, -45, -78, -59, 8, 17, -13, -32, 30, 14, -41, 2, 20, -18, 46, 36, 5, -17, -18, 0, 41, 12, -24, -19, 36, 1, -26, 12, 15, -22, -7, -26, 21, -15, 42, 1, -23, -15, 5, -35, -23, 28, 5, 19, -11, -37, 12, -8, 15, 0, 48, -17, 12, -23, 39, 0, 5, -18, -2, 46, 7, 1, -21, -4, -31, 13, 42, 32, -6, -15, -24, -52, -51, -13, 10, 14, 37, -28, -12, 42, 21, -24, 9, 55, -36, -27, 38, 12, -47, 7, 39, -11, -43, 44, 4, 7, -26, -7, -29, 32, 14, 8, -46, -47, 14, -27, 6, 0, -6, 43, -22, -3, 55, -21, -27, 39, -1, 10, -38, -43, 24, -4, 0, -9, -38, -7, 81, -13, 13, 14, -3, -45, 5, 12, 0, -29, 32, 42, 51, -32, 12, 20, -11, -7, -12, -56, 4, -4, 30, 34, 18, -51, -2, -39, -38, 3, 5, 21, 22, 48, 28, -58, -44, 15, -22, -3, -1, 30, 22, -42, -5, -8, 63, 57, 10, -23, -1, -63, 0, 25, -7, 7, 11, -46, -11, 49, 5, -15, -19, -35, 40, 28, 18, 17, -3, 2, -34, -65, -6, 24, -12, -1, 5, 39, -7, -20, -41, -25, 28, 3, -7, -8, -38, 1, -26, 13, -19, -11, -2, 4, -13, 6, -26, 24, -30, -10, 38, -10, 24, 24, -32, -14, 34, -2, 38, -13, -3, 20, -44, -21, -5, 28, 4, 57, 34, 5, -10, 2, 24, -54, -75, -4, 29, 20, -38, 34, 58, 10, -51, 14, 23, 8, -24, 25, -7, 36, -3, -12, -35, -8, -28, -7, -20, 20, 43, 5, -60, 20, 42, -27, 3, -25, -30, 47, 47, -36, 27, 0, 34, 22, 24, 10, -66, 12, -15, -47, 26, 42, -30, -6, 2, 3, 37, -25, -15, -25, 12, 23, 45, 31, -36, -25, -3, 47, 45, 32, -3, -5, -11, -24, -42, 37, 5, -36, -18, 23, -37, -53, 57, -10, -13, 14, -6, -23, -10, 21, -34, 3, 38, 20, 24, 38, -47, -73, 3, -18, 3, 21, 14, 45, 32, -25, 0, -49, -48, -7, 14, 30, -34, -57, 24, 1, -47, -30, -7, 17, 40, 39, 45, 13, -69, -49, -42, 52, -8, -41, 17, -17, -26, 51, 5, 18, 47, 58, -70, -19, 3, -44, -48, -18, 4, 44, 61, 21, -51, -38, 55, 70, -31, -10, 7, -6, -34, -3, -1, -12, 36, -20, -6, 9, 46, -40, 0, -18, 30, -1, -11, 14, -51, 11, -7, -13, 34, 72, 35, -15, -18, -34, -60, -27, 8, 36, 68, 8, -3, 13, -4, -10, -17, 0, 9, 6, 31, 7, -66, -20, -37, -20, 65, 21, 4, 46, 46, 11, -19, 0, -43, 30, -7, -14, 17, -37, -10, 31, 13, 39, 7, 8, -24, 21, -8, -41, 43, -29, 30, 39, 3, -48, 22, -11, -40, -30, -24, 55, 30, 29, 17, 44, 15, 1, 9, 12, -11, -42, -64, -44, 25, 25, 19, 54, -52, -5, 13, -35, -20, 30, -4, 39, 21, -48, -31, 26, -15, -4, 17, 21, 22, 9, -15, -4, -46, -31, -28, -21, 53, 41, 14, 5, 44, -46, -57, 54, 0, 14, 20, -32, -56, 63, 78, 38, -13, -1, -6, -64, 9, -19, -14, -48, -21, 38, -3, 0, 39, 44, -10, 7, -20, 12, -3, 1, -56, -48, 52, -2, -13, 25, 7, -59, 21, -20, -38, -45, 62, 4, -20, 59, 44, 24, -7, -41, 0, 14, -23, -8, -37, 10, -19, -23, -28, -18, -2, -8, 13, -11, 79, 39, -8, 17, 40, -48, -17, 48, 27, -1, -3, 27, -53, -57, 15, 71, 45, -75, -12, -15, -25, 39, 28, 44, 19, 17, -7, -55, -72, 21, 22, -28, -28, -27, 32, 36, 45, 5, 41, -21, 5, -17, -64, -44, 14, 39, 52, 14, -28, -31, -48, 30, -10, 10, 48, -6, -27, -29, 30, 0, -30, -22, -32, -8, 14, 5, -26, 42, -23, -47, 46, 0, -2, -8, 37, -2, 20, 31, 15, -5, -45, 12, -3, 0, -55, -31, -9, 72, 55, -20, -38, -39, 14, 58, -21, -15, -43, 13, -7, 10, -31, -39, 51, 54, 7, -2, 40, -18, -58, 5, -5, -12, -15, 28, 3, 30, -2, -43, -49, 13, -4, 21, 42, 55, -38, -47, -4, 4, -8, -22, -17, -3, -22, 20, 2, 28, -26, 8, 26, 36, -39, -68, -38, 49, 18, -5, 18, -22, -13, -35, -32, 60, 57, -18, -22, -4, 36, 20, -9, 37, 0, -11, 2, -21, -21, -27, -19, -49, 32, -6, -20, 59, 37, -12, 13, 27, -18, -7, -27, 28, -24, -31, 18, 62, -52, 18, -29, -40, 31, 32, -46, -8, 23, -4, 3, -42, -51, 65, 3, -38, 24, 24, -8, -36, 43, 0, -41, 32, 7, 31, -38, -44, 51, 71, 24, -34, -27, -68, -27, 26, -10, -24, 3, -15, 24, -4, -40, -43, 12, 14, 32, -7, 7, -17, 42, 25, 36, -71, 0, 48, -34, -6, -14, 38, 12, 54, -40, 21, 38, -8, -9, -34, -26, 40, -21, 39, -8, 19, 6, -25, -38, 4, 63, -30, -10, 28, -8, -63, 40, 0, 37, -27, 20, 15, 15, -53, 13, -30, 36, 55, -13, -40, 6, 25, -10, -9, -24, -11, 5, 26, 45, -17, 26, -10, 19, 20, 23, -71, -12, -21, 11, 40, -14, -42, -4, 15, 31, 4, -30, -46, 54, 61, 37, -4, -10, -27, -73, -43, 21, -10, -34, 29, 27, 26, 40, 14, 14, 20, -14, -46, 24, 21, -20, 19, -45, 4, -24, 40, -24, 48, 25, 7, -2, -56, -64, -11, 63, -30, 23, 18, -26, -1, 15, -5, -25, -12, 7, -1, 13, -27, -7, -4, -20, 35, 44, -22, -6, 27, 54, -40, 0, -7, -44, -6, 24, -47, -42, 0, -10, 44, -1, -4, -31, 12, 24, -27, -27, -24, 12, -20, -5, 31, 52, 40, -8, -1, -70, -40, 26, -13, 15, -1, 47, 20, 37, -18, -46, -18, -25, -24, 42, 8, 53, 30, 21, -27, -37, -8, 34, 23, -56, -9, -32, 49, 27, 22, 1, 11, -9, -55, -19, 36, 48, -18, -31, 37, 52, -4, -21, -26, -23, 21, 39, -21, -49, 10, 27, 8, -65, -17, -38, -13, -15, -3, -15, 36, 9, -28, 4, 63, -24, -56, -32, -3, 1, -10, 51, 46, -48, -3, 21, -17, 2, 57, -25, -27, 14, 21, 35, -8, -52, 39, -28, 25, 23, -10, 0, 13, 26, -29, 18, 5, -40, -65, -31, 11, 81, -12, 17, 21, -5, -52, 29, 42, -9, -38, -31, -1, 38, 0, 11, -44, -59, 42, -3, -32, 8, 25, 37, 0, -44, 12, 6, 2, 3, 7, 25, 24, -17, -31, 19, 25, -36, -6, 51, -25, -71, 27, -10, -34, -3, 31, -5, -8, 55, -27, -23, -2, -29, 53, -26, 14, 23, -7, 2, 0, 49, 38, -63, 3, -13, -7, -21, 3, 56, 26, 19, -4, 3, -8, -26, -73, 17, 1, -25, 0, -13, 47, -8, 30, 39, 1, -12, -37, -26, 38, 20, 27, -38, 29, -12, 8, 7, -12, 13, 20, -30, 24, -11, -47, 24, -8, -62, -40, 22, 1, 11, 5, 52, 23, -24, -48, -20, 26, 53, 32, 26, -65, -53, 9, -5, -21, 1, 54, 35, 21, -12, -14, 23, 20, 17, -29, -31, -34, 17, 59, 3, 19, -49, 12, 17, -35, -7, -7, -7, -21, -41, -21, 30, 3, 28, 75, 32, -1, 21, -12, -53, 18, 42, -32, 2, 25, 15, 6, -44, 4, 6, -27, -14, 41, 51, 25, -14, 0, -3, -37, -15, -6, 18, -39, -42, 29, 34, 39, 1, -40, 23, -31, 26, 44, -25, 2, 9, -18, -9, -23, -39, -6, -1, -23, 60, 4, 38, -29, 28, -21, -30, -21, -10, 0, -6, 12, 28, -13, -2, 27, 7, -41, 21, 26, -6, 14, 0, -21, -17, -21, -12, 18, -12, -44, -13, 71, 1, -12, -28, 18, 41, 21, -43, -39, 47, 40, 20, -34, 2, 31, -38, -42, -18, 22, 8, 51, -11, -57, 15, -3, 28, 25, 37, 18, 8, -37, -6, -19, 2, -2, 39, 53, -2, -3, -15, -26, -7, 0, -30, 1, 37, 54, 41, 26, -18, 15, 35, -59, -11, 31, -34, -52, 8, -10, 15, 34, 23, 31, -18, 21, -31, 7, 24, 23, -9, -46, -44, 24, 12, -23, -7, 40, 21, 7, -4, 8, 6, -34, -57, -42, 7, 88, 25, 13, 2, 19, -23, -72, 12, -1, 0, -18, -31, -3, 38, -25, -32, -31, 31, -28, 25, -15, -24, -13, 5, 25, 52, 22, -27, -29, -24, -22);

    signal memory_control : std_logic := '0';      -- A signal to decide when the memory is accessed
                                                   -- by the testbench or by the project

    constant SCENARIO_ADDRESS : integer := 1234;    -- This value may arbitrarily change

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);

                o_done : out std_logic;

                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,

                o_done => tb_done,

                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;

    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.

        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;

    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_rst <= '1';

        -- Wait some time for the component to reset...
        wait for 50 ns;

        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench

        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock


        for i in 0 to 16 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_config(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);
        end loop;

        for i in 0 to SCENARIO_LENGTH-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+17+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);
        end loop;

        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component

        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));

        tb_start <= '1';

        while tb_done /= '1' loop
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;

        tb_start <= '0';

        wait;

    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;

        wait until rising_edge(tb_start);

        while tb_done /= '1' loop
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH-1 loop
            assert RAM(SCENARIO_ADDRESS+17+SCENARIO_LENGTH+i) = std_logic_vector(to_unsigned(scenario_output(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(17+SCENARIO_LENGTH+i) & " expected= " & integer'image(scenario_output(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(SCENARIO_ADDRESS+17+SCENARIO_LENGTH+i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done == 0 before start goes to zero" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;

