-- TB EXAMPLE PFRL 2024-2025

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity tb_gen4_mod3 is
end tb_gen4_mod3;

architecture project_tb_arch of tb_gen4_mod3 is

    constant CLOCK_PERIOD : time := 20 ns;

    -- Signals to be connected to the component
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);

    -- Signals for the memory
    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    -- Memory
    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

    -- Scenario
    type scenario_config_type is array (0 to 16) of integer;
    constant SCENARIO_LENGTH : integer := 5000;
    constant SCENARIO_LENGTH_STL : std_logic_vector(15 downto 0) := std_logic_vector(to_unsigned(SCENARIO_LENGTH, 16));
    type scenario_type is array (0 to SCENARIO_LENGTH-1) of integer;

    signal scenario_config : scenario_config_type := (to_integer(unsigned(SCENARIO_LENGTH_STL(15 downto 8))),   -- K1
                                                      to_integer(unsigned(SCENARIO_LENGTH_STL(7 downto 0))),    -- K2
                                                      0,                                                        -- S
                                                      -1, 2, 4, -7, 8, -4, 0, 1, -9, 45, 0, -45, 9, -1           -- C1-C14
                                                      );
    signal scenario_input : scenario_type := (-31, 61, -25, -2, 57, -110, 21, -82, 62, 68, -35, 44, 68, -1, 78, -110, -96, -105, 70, 110, 65, -107, 126, -75, 74, -38, -82, 91, 85, -3, 70, -17, -26, 30, -99, 95, 103, 121, 4, -35, 82, 58, 25, 57, 112, 19, 42, 93, 28, -35, 7, -34, -75, -84, 93, -29, -62, -84, -108, -70, -72, 19, -125, -53, 107, -23, 88, 96, 81, -114, -42, -95, -101, -61, -63, -45, 90, -120, -48, -111, -4, 12, -60, -127, -32, -60, 126, -47, 75, -51, -110, 16, 29, -31, -52, -103, -18, -19, -95, -90, -1, -71, 45, 97, 96, 3, 114, 20, -27, -93, -64, -5, -54, 28, 39, 17, -10, 38, 77, 48, 26, -123, -71, -29, -66, -47, 58, 80, -74, -4, -99, 24, -109, 34, -70, 102, -6, 108, -112, -45, -1, -49, -14, 42, 108, -72, 65, -59, -30, -104, -48, -67, -47, 0, -55, -78, 6, -113, -126, -108, -72, 56, -19, 55, -80, -19, -109, 50, -3, -57, -95, 110, -4, 121, -122, -108, 22, -74, -23, 88, -32, 99, 62, -39, 72, -121, -102, -12, -69, 105, -105, 126, 120, -40, 72, 115, -106, 114, 107, 103, 120, 90, 69, -70, 106, -72, 3, 81, 13, 9, -121, -61, -83, -10, 71, 113, 80, -29, -50, 32, 17, -110, 45, -17, 56, -16, 22, -19, -122, 38, -14, 0, 99, -116, 127, -48, 123, -37, -93, -99, 78, -69, 60, 76, 115, -119, 11, -94, 20, 3, -101, 35, 79, 7, 124, -64, -91, -47, -92, -77, -110, -79, 57, 103, -125, 96, 28, -65, -76, 23, 49, -18, 91, -35, -58, 4, -50, -32, -126, -57, -113, 91, 28, 121, -100, 46, 103, -34, 126, 120, -51, 94, -79, -78, 4, 70, 30, -3, 60, -34, 11, 53, -15, -54, -26, 67, -43, 46, -33, -70, 1, 25, 44, -90, -23, -9, 73, 21, -20, 99, 120, 120, 73, 28, 35, -14, 108, -69, 66, 0, 24, 123, -71, -58, -91, 7, 67, -119, -39, 117, 115, 110, -43, -120, 79, 69, -1, 73, -81, 33, -31, -127, -40, -111, -7, 23, 103, 88, 55, 125, 70, 110, 3, -15, 57, -128, 87, -59, -114, 76, -13, 112, -106, 4, -24, 40, -70, -37, -79, 28, 97, -96, 24, 55, 66, -1, -104, 66, -57, 114, -73, 45, 48, -87, -5, 6, 14, -31, 127, 48, -89, -16, 33, 17, 24, -42, -30, 110, -40, 76, -55, -18, 55, -108, 4, -120, 75, -29, 88, -71, 48, 81, 69, -28, 3, 24, 57, -127, 88, -40, -5, 56, 37, -61, -3, 110, 113, -1, 126, 34, -3, 59, 99, 44, 34, -24, -114, 117, 37, 21, 51, -91, 67, 90, 118, 67, -56, 52, -56, 86, -52, 127, -63, 60, 38, 10, 84, 126, -65, -90, -86, 47, -27, 40, -69, -43, 108, -30, 29, 13, -43, -30, 125, 22, 115, 115, 11, 86, -8, 118, -125, 67, -74, -20, 57, 42, 57, -99, -99, 115, -104, -31, -10, -24, 114, 92, 45, -89, 0, 92, -13, 29, 77, 123, -120, -6, 85, -81, 24, -112, 116, 121, 106, -24, 61, 36, 122, 15, -65, 119, -122, -22, 31, 44, 76, -67, 102, 97, -14, -60, 107, 19, -33, -46, -46, -24, -33, 116, -18, 119, 60, -30, -117, 115, 118, -76, 14, 71, -2, -16, 24, -85, -84, 120, 105, 66, -41, -72, 94, 30, 106, -56, -73, -40, 115, 120, 94, 68, -22, -23, 43, 35, 57, 111, 38, -109, 119, 8, -35, 9, -104, 32, -80, -119, 32, 99, -103, 30, -114, 54, 27, -40, -71, -83, 96, 125, -94, -13, -3, 17, -16, 110, 122, -21, 27, -4, 110, -74, 91, 29, -119, -3, -57, 0, 16, -95, -6, -22, -90, -109, 117, 43, -27, 23, -16, 48, -80, 89, -65, 66, -108, 113, -110, -114, 48, 59, -77, 8, -91, 92, 84, 110, -64, -44, 34, 81, -15, 126, 72, 65, -77, 30, 98, -1, -72, 37, -106, 63, -93, -42, -88, 11, -61, -97, -122, -126, -31, 95, 67, -62, 59, 37, -120, 78, 78, -82, -114, 11, -103, -50, 14, -39, 75, -46, 100, 24, 78, 68, -35, -25, 9, -23, -70, -40, 14, -13, -9, 72, -56, 97, 97, 58, 54, -117, -18, 73, 117, -22, 1, 102, -23, -44, -37, 113, -107, 118, 75, 122, -49, 90, 122, 92, -3, -42, -48, 19, 2, 99, -52, 2, 38, 104, -43, -115, -81, -28, -112, -58, -107, 118, 114, 94, 72, 28, -22, 24, -24, 44, -99, -28, 107, -125, 47, 76, -25, -51, -77, -128, 81, -17, -59, 33, 41, 19, -108, -63, -102, -50, 112, -46, 64, -19, -112, -33, -46, 38, 89, -58, -21, -14, 122, -87, 6, -117, -6, 126, -2, 81, 34, -50, -35, 55, -32, -126, -61, 52, -87, -24, 18, 82, -46, 92, 96, 32, 30, -84, -42, 59, -124, 125, 67, 110, 59, 117, 17, -101, -24, 109, 109, -123, 95, -77, -89, 81, -65, 10, 127, 28, 126, 8, 88, 78, 45, 103, 73, -40, 47, 48, -124, -91, -81, -64, -94, -12, 109, -108, 0, -54, -118, -74, -127, 102, -100, 52, -25, 27, -115, -58, -55, -45, 87, -107, 81, -7, 60, -5, -64, -104, 0, 1, -42, 2, 119, 107, 127, -82, 47, -47, -92, 70, -4, -82, -53, -102, -84, -78, 3, -24, 10, 39, 26, 96, -53, 73, 67, -39, 89, 9, -48, -67, 84, 126, -96, 81, 25, 115, 114, -126, -98, -55, -87, 107, -85, 61, 98, -7, -15, 14, 26, 87, -89, -104, -30, -114, 42, -36, -4, 48, 2, -92, 108, -27, -102, -105, 8, -52, -10, -44, -127, 36, 67, -42, 85, 30, 70, -60, -91, 45, 126, -64, 84, 103, -14, -4, 46, 53, -112, -56, 56, -29, 78, -50, -46, -105, 115, 50, 26, -37, 43, 52, 78, 74, -72, 2, -88, -127, 117, 78, -14, -80, 94, -72, 27, -33, -19, -33, -62, 30, -109, -5, -63, 106, -50, -87, 111, 62, 39, -70, -113, -9, -59, -100, 19, 125, 33, 67, 4, 18, 102, 116, -15, 34, 56, -120, -78, -44, -41, 0, 15, -60, -127, -16, 44, -57, -11, 103, 94, -79, -113, -64, -71, -71, -121, 42, 67, 55, -100, 68, -104, -34, -41, -12, 17, -30, -32, 64, -71, -85, -77, 69, -100, -81, -67, 86, 16, -28, -1, 63, -1, 19, 56, -6, 89, 60, 87, -53, 125, 0, -26, -105, -79, -99, 42, -96, 125, 74, 70, -52, 40, 69, -113, 57, 127, -45, 16, -67, 25, 44, 70, -111, -127, 121, 7, 101, -29, 46, 36, 122, 32, -61, -61, 14, -36, -25, -71, -47, 62, 9, -85, 116, -26, 126, -10, -98, 31, 90, 27, 48, 35, 41, 79, -47, 126, 83, -39, 68, -107, -125, 58, -31, -123, -54, -98, 85, -48, -111, -86, 12, -85, -39, -41, -58, 44, 6, -20, 65, -30, -36, -93, 3, -119, 10, -15, -32, 118, -93, 48, -50, 75, -68, -93, 107, 123, 119, 7, -100, 109, 73, -4, -95, -47, -25, 80, 58, -2, 121, -3, 86, 115, 85, -73, 121, -38, -50, 43, 34, 73, 55, 4, 52, 111, -99, -19, 111, -7, -1, 124, 4, 60, 74, -69, 64, 39, -40, 104, -50, -10, 74, 76, -33, 126, -34, 26, -29, -91, -62, 82, -44, -117, 38, 46, 53, 107, -83, -57, -11, 19, -50, 80, -5, -52, 72, -64, -128, 70, -18, -126, -44, 69, 32, 112, 52, 86, 49, -51, 81, -121, 106, -15, -108, -16, -74, -67, 117, 114, -6, 64, 101, 30, -63, 77, 53, 41, 124, -10, 12, 100, 37, -74, 46, 48, -30, 108, -8, 26, 90, 85, -45, -48, -55, -17, 81, 23, -29, -18, 28, 126, -51, 60, -118, 127, -62, 95, -83, -19, -71, -75, 23, 15, -67, -127, -99, -24, -103, 77, -43, -44, -33, 81, 24, -124, -7, 118, 39, 81, 38, -72, 75, 28, 51, 13, -55, -70, 66, -74, 122, -57, 11, -31, 52, -29, 62, 98, -67, 58, 104, -84, -128, 116, -48, -28, -4, -43, -4, 64, -56, 18, -65, -127, 115, 120, 0, -122, 99, 65, 43, -62, 49, -61, 48, 107, 89, 93, 114, 28, -21, 64, 95, -22, -39, -86, -52, -1, 122, -25, -59, 17, -2, 45, 74, -89, -94, -116, -82, -127, -96, -75, -103, -120, 7, 10, -20, 85, -11, -9, 75, -52, -122, 100, -48, -68, 54, 32, 87, 125, -40, -33, 36, -80, -120, -4, -58, -107, -93, 125, -50, 25, -78, 4, -82, -5, -11, -52, -27, 92, 90, 84, -22, -71, 13, -126, 4, 37, -82, -119, -45, -28, -32, 100, -81, 74, -33, 62, -94, -40, 72, -41, 60, 29, -120, 47, -15, 89, 24, 102, 126, -21, -80, -84, 87, 22, -33, -108, -13, 105, -29, 39, -100, 88, 62, -101, -113, 90, 75, -109, -41, -66, -66, 36, 52, 80, 38, 124, -121, -5, 19, 114, -98, -68, 121, -79, 49, -107, 59, -64, -29, -66, 7, 75, -18, 53, 57, -41, 115, 71, 26, -16, 37, -63, -9, 80, 14, 103, 78, -22, -4, -6, 114, 86, 25, 82, 51, -128, -92, 56, 60, -9, -27, 95, -36, -74, -64, 98, -124, -23, 86, 72, 74, 97, 5, 9, 34, 11, 1, -39, 95, -75, -62, -80, -102, 77, 79, 68, 92, -64, -63, 35, 89, 30, -27, 127, -52, -25, 118, 40, 77, -23, -11, 54, 127, -74, -62, -32, 27, 113, 1, -48, 59, 36, -47, -14, 66, -25, -127, 51, -68, -60, -106, -24, -24, -59, 121, -77, -49, -103, 61, 90, 22, -76, 65, 18, 123, -6, -41, 105, 37, -89, -13, -84, 21, -27, 44, -82, -105, 87, 27, 46, -55, -124, -81, 30, -8, 20, 26, 79, -33, -2, -96, 14, 111, -113, 78, 33, 83, 99, 1, 25, 119, -29, -21, -66, 86, 0, -22, -125, -117, -16, -12, -72, 77, 2, 44, -89, -73, -55, 96, -17, -59, -108, 30, -85, 84, 85, -21, 62, -72, -49, -92, 24, -126, 127, 69, -21, 31, 80, -104, 80, 8, -27, -66, 125, -25, 125, 54, 22, 99, -18, 36, 40, -37, 1, 29, 70, 118, 65, -58, -65, 108, 69, -83, 86, 113, -95, -13, 89, -128, -61, 43, 65, -101, 89, 64, 111, 87, 80, -18, -96, 14, -25, -68, -76, -77, -95, 11, 25, -34, -13, -13, 15, 49, -13, 5, 68, 40, -47, 79, 46, 1, -20, 44, -124, -32, 48, 4, 14, 30, 119, 6, 55, 24, 27, 94, -4, -87, 108, -68, 81, 112, -15, 64, -42, -57, -2, -92, -110, -30, -92, -83, -93, -118, -44, -49, -28, -126, 20, 71, 27, 93, 61, 85, 45, -52, 111, 103, -47, 19, -21, -87, 100, 90, 17, -55, -33, 73, 77, -9, -19, 2, 65, 76, 69, -74, 35, -11, -115, 1, 5, 48, 75, -3, 24, -19, 71, -44, 126, -121, 87, -31, -97, -3, 12, 86, -60, -55, -128, -32, 67, -67, -71, 19, 101, -10, 76, -56, 79, 126, -62, -109, -91, -127, 90, -115, -80, 40, 34, -91, 70, -69, 10, 62, 53, -53, -18, -107, -67, 70, -7, 59, 108, 106, 31, 23, 40, 120, -88, -13, 115, 126, -98, -114, 80, -66, -112, 43, -96, -107, 91, 100, -94, -55, 18, -65, -5, 11, -39, -10, -52, -78, -71, -126, -15, 36, -106, -110, 100, 122, -103, -126, -121, -81, 4, 21, -37, -90, -91, 16, 62, -83, 61, -111, 99, 25, -36, -53, -31, -59, 93, 89, -50, -109, -9, 117, 49, 111, 7, -18, -71, -52, 64, -7, -108, 0, 16, 74, -12, 77, -52, -91, 10, 83, -40, 123, -15, -88, 22, 44, -31, -75, 5, -112, 75, -37, -128, 99, -73, 26, 27, 92, -69, -121, -18, 91, -82, -94, 59, -104, 10, 5, -10, 19, 30, 64, 67, 99, 81, -98, -128, -19, 98, 39, -61, -37, 25, -81, 17, 116, -17, 105, -82, -91, 39, -6, 120, -120, -7, 120, -45, 9, 69, -104, 60, 5, -17, 32, 58, 4, 54, -9, 32, -10, 29, 105, 29, -15, 76, 56, 81, 86, -45, -67, -114, -73, -80, 86, 79, -23, 96, 53, 114, 95, 56, 72, -86, 106, 20, -104, 115, 46, -128, -51, -101, -59, 72, -67, 50, 121, 57, -117, 95, -16, -13, 122, -39, 66, 44, -117, -62, 85, 30, -65, 56, 59, -124, -128, -16, 78, -6, 26, 112, 80, -83, 45, -116, 21, 25, -98, 14, 67, 77, -101, -82, -120, 123, 1, -111, -9, -23, 80, 56, -27, -59, -37, 25, -83, -43, -67, 104, 82, -75, 79, 38, -122, 13, -71, -47, -25, -93, 49, 35, -92, 57, 74, -87, 5, -113, -91, 43, 83, 29, 127, 121, -53, 83, -76, 104, 68, -69, 66, 43, 60, -28, 50, 105, -1, 30, 82, -23, 109, 107, 95, -97, -117, -51, 63, 126, 121, 17, 96, -49, -2, 95, 101, 89, -95, -13, -24, 98, -17, -67, -115, 75, 89, -23, -89, 26, -21, 45, -112, -77, -76, -13, -69, 110, -3, -38, -113, 95, 77, 3, -60, 127, -25, 73, 50, 85, 110, -97, -80, -8, -127, -71, -30, -56, 27, 16, 89, 38, 59, 120, -6, 107, 47, 37, 25, 81, 89, -6, -62, 97, 119, -49, -1, 65, -71, 40, 8, 62, 94, 54, 16, -15, 31, -97, 80, 53, 50, -25, 60, -110, -20, 77, 41, -84, 110, 127, -18, -106, 33, 12, -12, 57, 39, 112, 42, -102, -116, 89, -62, -38, -55, 43, -51, -120, 93, -70, -70, 38, -80, -81, -116, 56, 104, -5, 62, -83, 77, -60, -18, -85, 53, 87, 24, 104, -20, -98, 110, 109, 43, 125, 26, -94, -77, 104, -75, 75, -86, 122, -32, -86, -28, 57, -81, 96, 24, -101, 44, -27, -90, 85, 62, -35, 67, 1, -128, -22, -14, 36, -118, 88, -99, -64, -126, -8, -93, 121, 125, 47, -57, -37, 7, -83, -9, 113, 123, 10, 5, -108, -36, -89, 79, -28, -109, 13, 122, 93, 107, 21, -39, 112, -80, -127, 67, 86, -93, 103, -128, -120, 76, -18, -55, 72, 29, 20, -101, 100, -127, -9, -77, -42, -14, -84, -19, -121, 79, -37, -120, 39, -75, -89, 64, 97, 31, 1, -73, 19, -59, -98, -50, -43, -100, 6, -60, 112, -107, -52, -6, 105, -127, -17, -21, -28, -11, 26, -87, -61, -20, -22, 112, -84, -78, 5, -27, -121, -90, 94, 44, 60, -119, -115, -28, -7, 113, 124, 32, -61, 85, 65, 47, -9, -66, -119, -97, -38, 8, 34, 70, 81, 68, 24, -29, 83, -22, 97, 77, -78, 79, 124, 117, -6, -58, 33, 81, 54, -65, 122, 35, -79, 97, -126, 24, -62, 14, -24, 91, -3, 69, -20, 22, 43, -24, -53, -116, 115, -51, -4, -60, -51, -123, 78, -104, -106, -116, -67, 69, -98, 19, 23, -24, 92, 122, -21, -33, -1, -17, 111, -31, 35, 84, 27, -84, -118, -18, 109, 22, 114, -42, 71, 77, 99, -22, 85, -43, -69, -95, 23, -93, -24, 25, 23, 78, 64, 16, 64, 78, 58, 117, 22, 8, -30, -60, 23, -66, -6, -52, -10, -39, -122, -82, -20, 93, 3, -94, 114, -118, -76, -69, 71, 16, -96, 105, 70, 51, -70, -122, 36, -39, 42, -67, 104, 44, 103, -22, 118, -124, 105, 63, -117, -112, -119, 18, -64, 67, 59, 6, -61, 86, 35, -82, 17, -113, 50, -43, 33, 96, 1, 50, 43, 42, -123, -11, 99, -90, 76, 32, -121, -89, -64, -81, 27, -121, -37, 93, -33, -55, 56, 81, -35, -35, -86, 76, -84, -120, -39, 115, 121, 93, 21, 108, 67, 80, 100, -24, 75, 116, -124, -111, -101, -98, -47, 75, 63, -69, -101, 10, -84, 34, 123, -62, -115, -104, -115, 60, 60, -98, 113, -18, 86, -6, 5, 97, 105, -17, -62, 42, -1, -30, -105, -74, 119, 14, 88, -26, -117, 104, 45, -83, 76, 122, 49, 57, -56, 35, 48, -68, 24, -18, -113, -31, -74, -94, -80, 13, 19, -38, -45, 117, -53, 2, 5, 13, -23, -14, 72, 106, -50, -9, 120, 28, 28, 79, -32, 44, 92, -57, 116, 127, 99, -18, -57, -62, 68, -107, -91, 71, -72, -65, -91, -59, -28, -25, -57, 27, -38, 71, 40, -72, -75, 40, 56, -29, -6, 102, -73, -23, -20, 116, 70, 102, -60, -74, -52, 80, 66, 34, -105, -124, 26, 77, 2, 71, 18, -97, -75, 68, 116, 105, -30, -38, 51, 91, -7, -10, 55, 3, -59, -79, -6, 37, 117, 85, -119, 17, -121, 115, -126, 71, -37, -37, 39, -22, -115, 46, 18, 71, -61, -114, -91, 70, 56, 126, 8, -58, 22, 8, -5, -32, -3, -111, 33, -29, 81, 16, -16, 126, 16, -125, 66, -69, 18, 22, 107, 13, 3, 1, 48, 3, 42, 45, 106, -1, 40, 18, -51, 67, 35, -93, 15, -124, 101, 55, -27, 23, -79, -127, 111, -51, -125, -4, -27, -116, 32, 76, -58, -66, 69, 51, -52, 36, 14, -58, 34, -23, 47, -77, -96, 8, -16, -47, -29, 102, -106, -66, 100, 30, 8, -114, 67, -73, 32, 60, -86, -128, 25, 45, 29, -24, -46, -36, 61, -6, -25, 112, 125, 78, -79, 28, 79, -8, -74, -30, -73, 109, -13, -8, -82, 16, -3, 69, 57, 28, 29, -43, -85, 84, -103, -5, 38, 36, 1, -126, 56, -60, -14, 58, -20, 78, 15, -30, -44, 1, 100, -65, -119, 61, -16, 73, 71, 2, -6, 28, -19, -75, 99, -7, 89, 32, -14, 72, 68, 123, -65, 27, 73, 92, -90, 104, -100, -14, 25, 85, 27, -49, -86, 43, -127, -109, 107, -70, -37, 3, 26, 105, -30, 68, 10, 42, -15, 77, -84, 124, -32, -16, -113, -63, -119, 18, 45, 14, -114, 2, -108, 32, 6, 92, -103, 42, 65, 15, 14, -70, 15, 21, -83, -9, -119, -64, -55, -92, -78, 22, -17, 56, 122, -3, -22, -13, -32, -98, 70, -55, 115, 30, -86, 102, -51, -87, 60, -21, -87, 62, 94, -17, 109, 112, -92, -112, -28, 120, -9, -21, -91, -125, -122, -78, 39, 59, 86, 3, 61, -119, -26, 102, -117, -39, -61, -55, -37, -46, -68, -111, 5, -112, 117, -32, -103, -75, -125, -54, 15, 108, -22, 98, 84, 87, 9, -2, 111, -107, -101, -23, -33, -75, 16, 12, -91, 107, 26, -42, -93, 6, 70, 115, -121, -26, 104, -40, 15, 36, -114, 63, -41, -60, -120, 48, -101, -57, 62, -96, -10, 19, -40, -122, 43, -87, 77, 104, 63, -56, -8, 9, 30, -23, 108, -20, -111, 103, 96, 76, -127, -41, -56, -66, 51, -45, 97, 37, 118, -93, 49, 88, -22, 52, -34, 0, -35, 107, 56, 79, 38, 37, 48, -7, -7, 9, 81, -87, 33, -92, -12, -99, 4, 7, 122, -41, -83, 39, -26, 41, -17, -88, 20, 72, -57, -121, -1, -115, 39, -66, -81, 66, -57, 38, 24, -113, 2, -11, 117, 75, 119, 113, 29, 123, 93, 103, 39, 80, -20, 48, -71, -85, -105, 94, 49, -11, -110, -32, 95, -80, -89, 106, -97, 94, -50, 31, 46, -64, 81, 115, -71, 43, 122, 62, 102, -23, -69, -62, 58, 23, -42, 98, 41, 110, 62, 126, 95, 56, -117, -52, 4, -25, 73, 108, 112, 111, 58, 113, 115, 94, -65, -55, 6, -122, -102, 85, 117, -50, 67, 66, 33, 77, -3, 62, 29, 39, 121, 125, 76, -123, 35, 27, 60, 87, 106, 51, -75, 102, 62, 66, 66, 56, -72, 59, 45, -70, 4, -106, 46, -65, 90, 36, -116, 114, -48, 12, -31, 45, -123, 120, -30, 120, 31, 97, 34, 101, 20, 34, -21, 56, -73, -54, -10, 75, -75, 43, 2, 8, 4, 110, 11, 36, -94, 39, 90, -53, 36, 9, -76, 48, 24, -125, -127, 59, 110, 42, -126, -25, 20, -76, 31, 16, 105, -113, -111, -75, -125, -34, -76, 125, 6, 50, -118, 93, -11, 119, -40, -109, -34, 69, 124, -23, 85, -116, -20, 89, 24, 28, 86, -24, -34, 9, 22, -90, -82, 71, 45, 70, 20, -36, 41, 65, -9, -80, -88, 62, 116, 66, 60, 67, -59, 91, 104, -107, -91, 36, -12, 69, -69, 114, -123, -21, -121, -122, -115, -67, 71, 19, -63, -44, -13, 27, -55, -43, -117, -22, -78, 93, -1, -122, 19, -31, -89, -10, -49, -47, -5, -84, 42, 52, -27, 13, -117, -45, 65, -104, 97, 46, 55, 80, -108, -36, -73, 42, 116, -19, 41, 117, 10, 17, -71, 31, 126, 97, 4, 29, -48, -96, -56, 107, 105, -58, -29, -48, -80, 113, -58, 61, -94, 108, 79, -82, -75, 118, 58, 44, 94, 53, -20, -34, 37, -120, -36, 21, 82, 98, 11, 32, -101, -87, -121, -67, 103, -82, 92, 92, 6, 95, -9, -43, 117, -125, -65, -86, 50, -68, 45, -2, -125, -15, -70, 89, -63, -118, 44, -33, -45, 34, -57, 17, -36, 21, -90, -102, -106, -47, -95, -123, 64, 98, 14, 15, 31, -41, 41, 67, -15, 30, 111, -62, -120, -7, -117, -115, 111, -34, -89, 57, 98, 79, -27, -89, -108, -17, 122, 50, -58, 71, -58, -99, 15, 38, 52, -95, -65, 33, -65, 3, 112, -6, 97, -93, 112, 72, -94, -82, -46, 83, -88, -120, 96, -116, -20, 76, 10, 110, -10, 5, 109, 34, 119, 55, 107, 6, -62, 91, -24, -62, 68, -46, 91, -58, 101, 93, 12, -31, 114, -42, 96, 33, -46, -59, -75, -111, -2, -94, -56, 64, 85, -113, -29, 102, 99, -110, -63, -98, -11, -49, 20, 98, 59, -115, -87, 15, 80, -14, 13, 123, -3, 53, -119, -46, 50, -85, 124, 92, -119, -43, 0, -121, 57, -62, -122, 55, -34, 60, 3, 24, -72, 124, -36, -124, 38, -103, -95, 119, -101, 94, 108, 88, 2, 37, 126, 58, -42, 9, -15, -104, 41, 91, -45, -32, 6, -110, 18, -1, 90, 25, -99, 30, 10, 88, 43, -78, -14, 92, 122, -74, -121, -116, 123, -32, -25, -48, 12, 5, -118, -49, 29, -118, 38, -100, -77, -34, -99, -79, 7, 52, 38, -26, -49, 73, 124, -71, 119, 68, -13, -62, -85, 28, -115, 21, 88, -25, 44, -49, -81, -3, -116, -103, 3, 7, 83, 103, 35, -95, 109, 15, -61, -68, -90, 69, 110, 118, -16, -77, 7, -34, -25, -3, -12, -83, 84, -63, 9, 121, -118, 12, -6, -70, 95, -39, 100, 65, 79, -58, 35, 82, -109, -9, 18, 89, 63, -108, -105, 88, -66, 45, -70, -35, 49, 110, -103, 76, -82, 73, -86, -107, 7, 88, -6, -55, -47, 108, -83, -8, 106, -90, 54, 35, -123, 106, -15, -101, -43, 5, -110, 118, -33, -16, -113, -119, 12, -44, -118, 73, 59, 62, -8, 95, 95, -98, 33, 103, -58, 51, -14, 4, 121, -92, -126, -94, -88, -3, 62, 16, 70, 105, 72, 40, -72, -43, -7, 109, -94, 110, 108, 19, 103, -35, -120, 67, 35, 37, 126, 108, -42, 26, 69, -48, 80, -126, 104, -1, -39, 118, 84, 91, -103, -99, -78, 42, -101, 38, 75, 76, 114, 88, -91, 43, 122, -31, 90, 69, 121, 37, 117, 62, -20, 3, 58, -123, -25, 7, -43, -117, -84, -115, 12, 111, -95, 76, -101, 45, -112, 86, 127, 85, 35, -11, -16, 114, 17, 17, -29, 34, 20, -79, 121, -113, -44, -18, 23, 66, -69, 9, 75, -55, 96, 121, 71, -121, -11, -85, -67, 108, -12, -25, -102, 93, -39, 124, 98, -78, -123, -64, 98, -31, -127, -113, 55, -46, 91, -101, -32, -106, 40, -56, 24, 77, -76, 85, 68, -27, -102, -3, 103, -95, 117, -3, 5, 90, -82, 56, 23, -125, 17, 16, -69, -24, 52, -71, 73, -95, 104, 82, 76, 26, -64, -8, 87, 56, -86, 62, -115, 67, -112, -68, 47, 118, 2, 4, -119, 108, 113, -12, 119, -50, -13, -102, 70, 37, -52, -111, -11, -122, 45, 91, -28, -89, 59, -86, -40, 126, -119, -50, 13, -115, -64, 34, 68, -87, 24, 21, -122, 64, 81, -104, -28, -44, 74, 78, -53, 23, 32, 61, 84, -88, -69, -32, 90, -116, -117, -37, -65, -35, -46, 97, -50, 84, 49, 54, 36, 113, 122, -40, -113, 0, 116, 117, 117, -64, 7, -4, 25, 10, -106, 80, -79, -119, 83, 28, 55, -41, 66, 97, -53, -90, -66, 116, -52, -39, -64, 42, -57, 85, 62, 79, 14, -34, -22, 7, -36, -6, -61, -64, 120, 12, -93, -69, 87, 32, 11, 10, -103, 106, 46, 69, -83, -55, 68, 126, 91, 116, 65, -76, 82, 45, -91, 119, 100, -61, 82, -101, -77, -52, 15, -78, -61, -34, 123, 22, -89, 43, -125, -117, -4, 114, -51, -123, 112, -15, -95, 106, -31, 25, 121, 102, 115, 4, -52, -80, -42, 12, -25, 89, 51, 9, 67, 44, 127, -123, 117, -75, -115, -89, 71, -93, -106, -76, -111, 11, -12, 51, 7, 48, 37, -128, 12, -3, -25, 36, 2, 79, -106, -110, -63, 121, -13, -25, 12, 27, -117, -76, 100, -127, 40, -92, -37, 21, 68, -102, 123, -76, -12, 28, 45, 72, 81, 33, 97, 49, -67, -52, -55, -117, 75, 124, -57, -80, 44, 91, -35, 122, 55, -42, -59, 33, -104, 99, 29, -25, -50, 47, -93, -46, 105, 97, 45, -128, -119, 125, -3, 46, 115, -8, 105, -121, -52, -4, 38, -25, -59, 27, -86, -76, -67, 125, 103, -47, 60, 106, -85, -64, 10, 24, -117, -66, -43, -22, -120, 76, 41, -127, 116, -107, -99, 86, 54, 63, 88, -115, 7, -123, 15, -51, -113, 64, -72, 41, 107, -108, 103, 5, -88, 94, -28, -125, -4, 84, -7, -26, 4, 15, -25, 6, -76, -82, -52, -80, -27, 58, -127, -89, -45, -22, -52, 40, 8, -4, 111, -36, 123, 108, -76, -58, 106, -28, 41, -107, 32, 8, 46, -11, 104, -87, 23, -19, 110, -66, 59, 32, 110, -14, -48, 110, -120, 34, -40, -92, 58, 104, -44, 99, 121, -84, 32, -90, 47, -39, -96, -46, 11, -125, 123, 66, -10, -7, -38, -78, 15, 83, -21, 61, -20, -34, -121, 73, 29, 54, -29, 78, 35, -90, 63, -103, 72, -126, -103, 32, 30, 108, 16, 26, -123, -71, 73, -61, 106, 52, -61, -120, -85, -98, 46, 51, 66, -101, -85, -1, -80, -102, 91, 4, -55, 110, 82, -120, -90, -97, -90, -86, 51, -111, -56, -87, 53, -31, -93, 86, -91, 6, 42, 83, -87, 11, -73, 75, -26, 3, -41, 87, -22, -111, -25, 5, 8, -33, 8, -55, 39, 14, 34, 107, -20, -13, -73, -26, 90, -81, 75, -102, 96, -7, -122, -72, 126, -17, 46, -92, -106, -127, 76, -17, -32, -25, -54, 62, 3, -126, -2, 29, 25, -32, 40, 10, -100, 67, 31, -86, 51, -42, 107, 125, 44, -108, -64, 45, 53, 33, 72, 111, -52, -91, 6, 17, -29, -35, 33, -120, -27, -125, 107, -52, -119, -127, 127, -106, 31, 4, 114, 95, 79, 23, -33, 63, 112, 21, -101, 124, -29, 25, 103, -78, 70, 44, 103, -73, 12, -40, -110, 103, -34, -58, 68, -98, -48, -124, -126, -29, -27, 125, 83, 55, 36, 12, 69, 110, 112, -110, -93, 21, -73, -34, -90, 10, 6, -117, 76, -58, 10, -2, 57, 55, -24, 93, -115, -128, -4, -1, -95, 79, 17, 63, -111, 77, -63, 73, -63, 32, 36, -73, 112, 80, 104, -80, -92, 43, -98, 74, -100, 72, 102, -25, -18, 121, -54, 75, -10, 24, 109, -57, 5, -54, -79, 54, -25, -83, -17, 35, -35, 87, -95, -126, 62, 89, 125, -117, 117, 105, 41, 116, -30, 64, 48, -80, -128, -42, -73, 70, 60, 50, -50, -60, -81, 105, 67, 59, 35, 14, 94, 37, -4, -60, 117, 83, 33, -107, 44, -121, 74, 117, -63, 110, 43, 52, 90, -104, -40, -43, 36, 77, 2, -24, 93, 42, -113, -53, 80, -16, 32, -6, -29, 88, -16, 96, 127, -121, 101, -49, 30, -106, 123, 60, 64, -72, 14, -92, 57, -110, 54, 123, 123, -56, -3, -35, 67, -47, -41, 9, 53, 73, -31, 109, 88, -33, 40, 67, 15, 3, 99, -51, -49, 100, 75, -67, 62, -69, 48, -53, -13, 22, 111, -89, -85, 16, -2, -94, 34, 11, 47, 110, -89, -75, -100, -17, -83, 37, 0, -65, -90, 12, 18, -14, -44, -35, -102, 71, 66, 70, -16, 21, -126, 35, 56, 81, 51, 108, 71, -122, 17, -77, 43, 52, -38, -20, -81, 22, 99, 74, -29, 44, 121, -21, 18, -51, -42, -27, -19, 66, 72, 107, 125, -103, 58, -124, -78, -38, 65, 7, 71, -120, -57, -69, -97, 1, -92, 66, -111, -58, 89, -128, -94, -110, -95, 113, 45, 21, 123, 47, -97, 4, -30, 20, -112, -52, -4, -112, -88, 126, 80, 90, 88, 99, -73, -48, 67, -101, -123, 107, -71, 49, -82, -42, 124, -94, 23, 74, 38, -68, -64, -24, 37, 98, 115, -9, -109, 3, 90, 101, -85, 35, 121, 91, -27, -14, -17, 92, 31, 85, 12, -78, -24, -54, -126, -74, -93, 61, -91, -117, -55, -79, 38, -125, 106, -90, -47, -112, -119, -57, 63, 70, 109, 113, 28, -61, -104, -26, 53, 84, 102, -23, 83, 90, -42, -62, 19, 4, 7, 72, -91, -118, -16, -81, -36, 100, -82, -31, -128, -110, 11, -18, 46, 31, -11, -89, -109, 38, -93, -65, -27, 9, 30, 15, 32, 69, -41, -74, 107, 12, -82, 90, -51, 57, 119, 15, -30, 125, -65, -89, 9, 11, -117, 8, -62, -86, 120, 76, 47, -59, 126, 56, 97, 86, -66, 1, -76, 124, -98, -32, -25, 45, 35, -61, -127, -122, 63, -24, 102, 66, 27, -115, 80, 38, 115, -80, -58, -30, 117, 46, 79, -112);

    signal scenario_output : scenario_type :=(65, -59, 8, 75, -116, 122, -113, 53, -2, -68, 58, 17, -55, 117, -73, 58, -58, 18, -38, 18, -101, 127, -128, 127, -43, -48, 76, -27, -55, 96, -28, 5, 71, -123, 91, -53, 32, -5, 3, 74, -27, -12, 17, 50, -42, 31, 50, -6, -2, 58, -7, -5, -52, 88, -92, 18, 21, -23, 1, -60, 53, -111, -2, 69, -128, 65, -3, 59, -59, 111, -28, -23, 0, -38, -58, 93, -128, 96, -68, 21, -12, -23, -33, 53, -113, 101, -128, 123, -33, -29, 58, -23, -31, 28, -36, 29, -12, -44, -12, 38, -106, 22, -16, 8, -50, 113, -26, 37, 0, 6, 15, -76, 23, -13, -6, -10, 16, 11, -8, 59, -43, 49, 6, -53, -32, 11, 16, -80, 108, -80, 95, -128, 98, -128, 102, -114, 127, -106, 69, 21, -58, -1, -15, 57, -118, 127, -70, 57, -43, 29, -38, -24, 13, -36, -28, 66, -69, 6, -10, -63, 27, -103, 78, -74, 85, -93, 75, -49, -5, -57, 108, -128, 127, -97, 29, 79, -109, -11, 59, -123, 88, 0, -55, 127, -90, 23, 44, -127, 122, -128, 127, 1, -95, 92, 74, -128, 127, -44, -12, 43, 17, 71, -70, 127, -119, 38, 39, -50, 64, -45, 60, -53, -21, -21, -8, 17, 0, 16, 47, 6, -93, 109, -88, 47, -47, 44, 17, -75, 96, -73, -31, 103, -128, 127, -128, 127, -58, 24, -28, 93, -128, 63, -31, 78, -113, 127, -95, 49, -5, -88, 58, -2, -86, 127, -66, 33, 49, -47, 7, -38, -47, 0, 31, -128, 127, -38, -22, 3, 24, -10, -73, 101, -53, 6, 54, -48, 39, -59, 52, -117, 74, -119, 107, -127, 97, 38, -123, 103, 28, -97, 127, -75, 13, 12, -3, -29, -13, 73, -54, 27, 31, -23, 0, -3, 52, -98, 81, -27, -17, 28, -26, 32, -68, 57, -37, 23, -27, -33, 54, -18, 13, 24, 23, 54, -43, 117, -128, 116, -49, -12, 101, -90, 75, -31, 3, 38, -116, 26, 32, -58, 50, 3, -24, 101, -45, -57, 111, -95, 101, -11, -53, 76, -93, 16, -55, 3, -11, -16, 71, -28, 79, -11, 16, 107, -128, 127, -81, -57, 114, -128, 121, -127, 106, -47, 45, -63, 49, -54, 7, 45, -128, 90, -13, 3, 16, -57, 127, -128, 127, -128, 81, 28, -79, 66, -17, 0, -68, 91, -18, -43, 65, 3, -34, 27, -18, -18, 92, -128, 122, -68, 18, 75, -118, 118, -128, 111, -128, 102, -109, 69, -5, 11, -23, 45, -1, 60, -128, 127, -107, 8, 27, 3, -42, 16, 22, 0, -70, 127, -29, 0, 38, 21, -18, 45, 32, -79, 127, -91, -3, 80, -97, 87, -38, 10, 33, -37, 127, -101, 113, -128, 127, -128, 96, -11, -32, 29, 64, -54, 59, -18, 48, -100, 65, -54, -13, 90, -116, 59, 12, -21, -26, 79, -112, 59, 32, -44, 109, -69, 127, -128, 127, -101, 11, 21, -42, 59, -42, -18, 127, -128, 63, 2, -73, 49, -28, 38, -33, 49, 42, -86, 29, 3, 81, -117, 90, 65, -128, 124, -128, 95, -53, 27, -36, 96, -39, 69, -15, -43, 127, -128, 73, -1, -39, 52, -101, 106, 0, -22, -16, 109, -58, 6, 27, -2, 0, -68, 86, -128, 101, -5, 18, -57, 103, -6, -102, 87, 32, -44, 7, 63, -47, -38, 68, -63, 21, 11, -13, 91, -98, 90, -47, 36, -22, 24, -42, 1, 54, 3, 21, 32, -31, -7, 45, 21, -86, 127, -79, -8, 80, -93, 103, -64, -48, 34, 27, -128, 127, -127, 85, -31, -17, 21, -53, 38, 17, -111, 102, -8, -1, -58, 45, 21, -58, 88, -39, 103, -128, 127, 0, -74, 109, -69, 6, 22, -78, 63, -8, -27, -65, 92, -79, -28, 68, -39, 69, -111, 127, -128, 127, -128, 127, -123, -7, 58, -17, -90, 107, -109, 74, -60, 58, -47, 45, 16, 12, -93, 100, -36, 64, -52, 64, 32, -34, -21, 116, -128, 127, -112, 57, -55, 48, -49, 0, 0, -43, -33, -2, -21, -71, 100, 18, -116, 116, 0, -54, 6, 92, -108, 6, 17, -91, 81, -116, 102, -69, 38, 34, -23, 34, 26, -10, -18, 2, 8, -37, -23, 68, -114, 86, -16, -11, 88, -65, 57, -8, 15, -59, 29, 86, -60, 28, -26, 112, -128, 127, -74, 73, -87, 98, 1, 11, 12, 38, 0, 24, -64, 78, -87, 50, -10, 52, -36, 15, 24, 18, -81, 37, -117, 63, -68, -5, 39, 32, 0, 55, -45, 78, -85, 12, 101, -128, 108, 6, -47, 37, 24, -87, 98, -92, -33, 48, -18, 24, -42, 66, -45, -48, 73, -128, 102, -7, -37, 60, -63, -6, 33, -75, 58, -39, 100, -128, 127, -87, 8, 48, -121, 81, 11, -13, 11, 54, -29, -31, 12, 49, -119, 33, -21, 34, -106, 85, -1, -21, 74, -31, 15, 79, -128, 127, -95, 33, -18, 85, 13, -18, 29, 17, 23, -128, 127, -97, -28, 116, -128, 12, 59, -102, 107, -65, 73, 8, -17, 57, 28, -42, 78, 43, -69, 59, -11, -13, -60, -23, 71, -128, 113, -12, -38, 42, -121, 127, -128, 112, -70, 69, -70, 49, -21, -64, 90, -128, 127, -91, 53, -5, 12, -22, 36, -28, -44, -12, 27, -45, 88, -87, 127, -32, -53, 92, -52, -24, 54, -34, -1, -45, 8, -58, -3, 3, -36, 78, -98, 92, 12, -76, 112, -29, 7, -26, 36, 34, -128, 127, -76, 33, 70, -73, 80, 24, -113, 113, -128, 76, 21, -48, 31, 22, -24, 73, -63, 24, 60, -119, 76, -88, -1, 27, -2, -80, 127, -74, 2, -3, 44, -86, 22, 2, -80, 57, -10, -102, 97, -53, 68, -24, -11, 31, 37, -128, 107, 23, -49, 36, 26, 39, -70, 33, 49, -113, 93, -60, 53, -81, 96, -81, 21, -16, 48, -23, 3, 50, -54, 108, -27, -80, 95, -66, -8, -29, 127, -128, 87, -37, 12, 2, -42, 75, -112, 78, -103, 102, -86, -38, 102, -71, 33, 6, -7, 60, -48, -58, 7, 16, -80, 66, -8, 2, 29, 28, -49, 66, 69, -75, 54, 0, -45, -7, 7, -11, -37, 29, 5, -85, 2, 31, 13, -34, 38, 34, -34, -5, -86, 38, -48, 23, -91, 127, -119, 55, -26, -16, 7, -28, -21, 75, -69, 24, -36, 81, -117, 34, -45, 45, -64, -8, 12, 34, -47, 13, 36, -58, 63, -32, 68, -91, 127, -65, 48, -6, 31, -70, 71, -128, 111, -69, 44, -42, 68, 53, -128, 90, 38, -107, 109, -54, 37, -27, 53, -52, -28, 124, -128, 91, -69, 68, -34, 58, -8, 6, 18, 39, -52, 21, -26, -23, 36, -27, -86, 127, -128, 124, -34, -31, 64, -1, -54, 37, 5, 0, 63, -97, 114, -6, -60, 127, -66, -23, 96, -70, -45, 65, -107, 90, -85, -3, 1, 39, -96, 26, -10, -54, 38, -38, -32, 71, -49, 42, -38, 76, -119, 64, -43, -66, 122, -128, 127, -96, 100, -65, -38, 71, -59, 24, 26, -45, 127, -44, 5, -2, 42, -47, 15, -22, -50, 113, -91, 58, 16, 39, -85, 127, -88, 2, 52, -48, 15, 10, -15, 24, 86, -103, 52, 70, -90, -3, 96, -90, 52, 57, -88, 102, -7, -71, 127, -96, 24, 28, 6, -81, 127, -101, 80, 5, -18, -18, 68, -71, -45, 74, -53, -32, 88, -71, 55, 8, 2, -81, 87, -44, -36, 109, -58, -53, 116, -63, -54, 26, 15, -90, 52, -34, 52, 33, -50, 127, -128, 127, -59, -42, 88, -54, -60, 49, -23, -60, 68, 34, 1, -38, 95, -37, -28, 91, -58, 27, 63, -5, -49, 86, -2, -78, 113, -76, 22, 29, 24, -27, 53, -2, -28, 28, -34, -1, 15, -16, 71, -118, 127, -128, 127, -128, 127, -101, 78, -22, -34, 26, -16, -13, -2, -2, 21, -128, 98, -95, 13, -23, 42, -7, -70, 48, 31, -91, 54, 33, -59, 107, -57, 24, 17, 0, -22, 92, -128, 127, -123, 76, -42, 54, -76, 36, 48, -102, 85, 55, -64, -28, 127, -128, 27, 29, -39, -3, 47, -87, 86, -17, -87, 91, -38, -11, -53, 127, -68, 23, -43, 112, -97, 36, 1, -27, 13, 57, 3, 1, 49, 29, -37, 55, -7, 0, -44, 55, -74, 8, 55, -48, 1, 53, -54, 58, -11, 7, -57, -10, -13, -36, -60, 23, -45, -63, 74, -57, 0, 80, -39, -58, 127, -114, -21, 64, -68, 3, 64, -52, 44, 75, -49, -24, 64, -52, -26, -58, 107, -128, 96, -60, 73, -74, 34, -12, -32, -22, 26, -37, 34, 5, 3, 97, -118, 54, 8, -54, -2, 26, -33, -70, 93, -128, 127, -95, 101, -81, 17, 63, -116, 69, 22, -97, 123, -100, 53, -65, 37, 52, -22, 44, -23, 68, -64, 15, -24, 11, 44, -113, 107, -109, 102, -2, -50, -10, 75, -18, -90, 96, -21, -47, 15, -44, 10, -37, 127, -122, 107, -39, 73, -101, 11, 127, -128, 127, -123, 123, -93, 39, -38, -1, 23, -79, 50, 26, -81, 102, -31, 11, 3, 73, -59, 12, 37, -81, 57, 15, -21, 53, -32, 44, -18, -22, 69, 49, -50, 24, 34, -39, -27, -13, 96, -63, 18, -27, 112, -128, 48, 21, -53, 0, 55, -17, 34, 29, -7, 18, -47, 111, -96, 52, 6, -78, 45, -59, -22, 79, -37, 24, 23, -2, -21, -39, 127, -102, 11, 80, -81, 69, -22, 18, 3, 68, -85, 60, 1, -32, 36, -44, -8, 71, -8, -33, 16, 49, -23, -65, 127, -100, 29, -39, 21, -26, -90, 127, -127, 74, -64, 39, -24, -7, -43, 102, -87, 79, -43, -13, 98, -21, -47, 98, -76, 50, -73, 64, -49, -38, 88, -95, 43, 1, -2, -1, 17, -74, 5, -16, 52, -53, 78, -63, 21, 69, -128, 127, -68, 8, 38, -31, 22, 90, -70, 66, -48, 81, -66, 43, -15, -6, 15, -32, -90, 85, -81, 69, -45, 34, -47, 59, -75, 28, -34, 87, -128, 66, -7, -68, 117, -58, 54, -52, 80, -128, 124, -57, -42, 48, 71, -128, 127, -52, 7, -52, 119, -128, 108, -29, -11, 96, -64, 55, 27, -37, 29, -8, -13, 24, 21, -2, -3, 75, -18, -97, 107, 38, -108, 66, 95, -128, 45, 13, 8, -128, 123, -66, 18, 2, 54, 18, -15, 78, -34, -15, 7, -1, -57, 15, -22, -43, 24, -11, -7, 21, -34, 6, 31, 1, -55, 88, -23, 0, 0, 88, -102, 44, 13, -58, 6, -16, 63, -69, 68, -2, -6, 64, -13, -53, 127, -128, 75, 26, -78, 114, -31, 5, 57, -48, -17, 42, -66, 0, -8, -50, 10, -50, 16, -96, 44, -17, -66, 50, -18, 39, 32, -57, 97, 8, -68, 97, 5, -78, 80, -34, -2, 10, 5, 26, -7, -24, 28, 0, 7, -11, 47, -63, 103, -1, -69, 66, -52, -13, 23, -34, 54, -37, 78, -113, 127, -128, 127, -55, -34, 53, -54, 50, -66, 69, -47, 2, 32, -91, 1, 7, 23, -95, 111, -92, 65, 50, -59, 47, 44, -107, 121, -128, 7, 37, -15, -101, 127, -113, 32, 5, 7, -36, 79, -45, -18, 48, -102, 17, 10, 13, -2, 34, 0, 97, -106, 49, 31, 28, -63, 13, 127, -106, -42, 116, -100, -48, 63, -6, -88, 58, 49, -85, 26, 3, -39, 34, -12, -6, 18, -70, 13, 12, -78, -33, 58, 2, -80, 71, 5, -42, -16, -22, -17, 0, -21, 6, 12, -119, 127, -128, 127, -53, -5, 18, 21, -73, 45, -2, -26, 3, 15, 21, -92, 78, -16, 50, 1, -17, 47, -33, -53, 64, -49, 24, -69, 101, -38, -8, 26, 22, -124, 127, -49, -22, 65, -3, -27, -13, 79, -128, 114, -59, -88, 127, -128, 59, -33, 63, -44, 0, 18, 45, -100, -6, 114, -128, 68, -22, -28, 10, -13, 6, -11, 24, 59, -24, 21, 8, 3, -36, -21, 29, 49, -95, 21, 48, -119, 127, -69, 5, 69, -109, 119, -128, 63, 76, -122, 47, 78, -128, 121, -47, -21, 22, 12, -38, 59, -34, 47, -27, 0, 44, -27, -11, 65, -32, 13, 54, -21, 59, -11, 13, -87, 32, -27, -75, 98, -50, 39, 10, 3, 93, -98, 127, -28, -96, 127, -23, -71, 107, -50, -42, 59, -128, 44, 21, 10, -92, 127, -90, -26, 111, -123, 88, 34, -65, 23, 49, -47, -59, 76, 29, -64, 21, 5, 0, -81, 6, 42, 22, -73, 127, -122, 71, 5, -95, 54, -16, 32, -58, 78, -92, 106, -86, -48, 86, -71, 24, -8, -7, 18, 1, 39, -75, 43, -75, 50, -8, -98, 127, 7, -92, 127, -71, 1, 18, -90, 57, -8, -97, 86, 18, -97, 123, -63, -21, 15, -27, -70, 59, 45, -85, 127, -128, 108, -2, -85, 108, -39, 33, -43, 39, 39, -57, 34, 59, -88, 80, -16, 64, -26, 43, -2, -24, -28, 12, -37, 127, -59, 28, 28, -24, 60, -59, 98, -55, 63, -54, 31, -49, 59, -24, -29, -11, 80, -75, 71, -75, 49, -29, 12, -111, 96, -75, 37, -65, 88, -47, -8, -39, 127, -128, 76, -23, 10, 81, -64, 54, 68, -97, 18, -2, -71, 22, -55, 34, -34, 8, 73, -80, 107, -24, 22, 1, 28, 27, -3, -26, 71, 16, -76, 59, 69, -106, 86, -49, 6, 16, -1, 24, 3, 74, -109, 98, -53, 18, -33, 114, -100, 38, 22, -12, -92, 103, 5, -27, -8, 93, -44, -38, 39, -44, 53, 17, -8, -13, 118, -128, 37, -32, 53, -42, -74, 127, -123, -6, 81, -80, 31, -66, 28, -12, -81, 113, -100, 127, -95, 60, -69, 37, -11, -64, 97, -17, -49, 102, -39, -54, 102, 7, -2, -1, 111, -128, 127, -128, 127, -76, -2, 21, 45, -128, 116, -22, -75, 118, -42, -73, 86, -29, -66, 97, 2, -59, 74, -49, 42, -128, 127, -127, 65, -59, 59, -128, 68, -33, 1, 7, 42, 42, -75, 0, 11, -3, -28, 92, -37, 70, -97, 80, -63, -47, 33, 1, -55, 50, 13, -23, 127, -85, -28, 79, -5, -128, 127, -119, -10, 98, -97, -43, 74, -48, 43, -88, 127, -128, 108, -55, -1, 15, -66, 63, -123, 113, -71, -63, 119, -87, -42, 42, -23, -28, 48, -27, 78, -39, -18, 21, -7, -74, 57, -118, 127, -128, 54, -24, 78, -128, 101, -17, -28, -8, 37, -58, 22, 3, -73, 97, -103, 27, 47, -18, -44, -27, 53, -93, 68, -44, 28, 18, -81, 8, 0, 5, -26, 100, -34, 12, 23, 26, -2, -5, -21, -33, -32, -2, 2, 17, 23, -23, 97, -98, 73, 26, -92, 97, -13, 18, 1, 12, 44, -2, 10, -80, 127, -32, -73, 127, -128, 127, -85, 38, -69, 68, -80, 78, -45, 32, 27, -17, 33, -85, 127, -128, 64, -16, 31, -97, 127, -127, 32, -13, -50, 59, -128, 71, -7, -68, 44, 28, -45, 44, 36, -59, 87, -101, 45, 33, 2, 1, 0, -2, 21, -111, 108, -91, 86, -16, 43, -60, 127, -44, 33, -29, 69, -108, 21, -3, -47, 21, 2, -16, 39, 10, -21, 71, -22, 49, 21, -22, 60, -78, 48, -44, 22, 1, -42, 7, -42, 23, -38, -73, 127, -128, 60, -44, 34, -32, -95, 117, -58, 33, 3, -22, 92, -111, 63, -109, 98, -78, 71, -79, 127, -128, 127, -1, -60, 69, -47, 44, -128, 47, -18, 1, -39, 91, -17, -59, 121, -121, 103, -101, 11, 36, -66, 53, 1, 58, -78, 50, 66, -128, 121, 2, -57, 53, 0, -73, 68, -119, 8, 57, -88, -10, 45, 7, -48, 59, -58, 109, -93, -6, -8, 3, -48, 15, -15, 87, -21, 18, 66, -59, 70, 80, -91, 80, 7, -47, -49, 6, -10, -29, 2, 78, -116, 15, 54, -75, 38, 33, -81, 31, -16, -128, 127, -127, 90, -42, 0, 37, 17, -17, 5, 74, -36, 17, -18, -36, 75, -128, 85, -3, -64, 127, -44, -90, 90, 0, -44, 79, -44, 65, 23, -76, 80, -2, -55, 65, -38, -21, -31, 5, -23, -28, -36, 111, -123, 59, 0, 3, -15, -13, 13, 34, -68, 28, 74, -69, 12, 74, -66, 47, 54, -118, 103, -17, 26, 10, 45, -18, 93, -109, -8, 98, -113, 36, -13, -8, -15, -15, -49, 49, -86, 53, 0, -27, 2, 32, -11, -47, 3, 93, -106, 65, -44, 44, -64, 79, -31, 47, -18, 26, -42, 34, -11, -6, 33, -22, -76, 68, 15, -24, 1, 18, -36, 21, -16, 28, 32, 13, -42, 16, 52, -13, 1, -5, 8, -45, 11, 37, -88, 127, -128, 127, -128, 127, -74, -12, 52, -16, -70, 90, -78, 52, -28, 15, -24, 31, -93, 54, -16, 0, 68, -22, 0, -10, 52, -93, 88, -101, 55, -33, -37, 106, -22, -73, 127, -128, 44, -42, 47, -43, 32, 3, 32, -37, 26, -18, 57, -52, 63, 22, -52, 73, 0, -71, 127, -128, 109, -50, -43, 91, -22, -70, 127, -111, -34, 78, -26, -92, 52, 7, -68, -1, 58, -18, -63, 75, 0, -53, 73, -65, 70, -47, -8, 47, -43, -24, -28, 100, -123, 12, 74, -78, 47, -74, 127, -128, 45, 34, -49, -16, 55, -49, -10, 1, 11, -18, 43, -49, -34, 53, -15, 36, -45, 81, 24, -28, -2, 55, -92, 95, -97, 52, -39, 53, -60, 18, -8, -1, 45, 1, -43, 127, -128, 55, -3, -15, 32, -81, 127, -108, 3, 42, -86, 73, -21, 7, 5, -12, 66, -66, -27, 108, -118, 33, 7, -15, 21, 38, -5, -60, 108, -118, 70, -10, -22, 57, -34, 85, -88, 80, 0, 45, -117, 127, -128, 58, -17, 10, -7, 11, -17, 108, -108, -32, 121, -128, 31, 8, -42, 57, -93, 97, -37, 43, -44, 101, -128, 127, -101, 70, -33, 50, -87, 24, -33, 6, -65, 114, -117, 63, -78, 81, -127, 96, -3, -33, 50, -42, 49, 10, -69, 90, -74, 27, -8, -43, -32, 24, -81, 0, 45, -48, 39, 32, 10, -75, 108, -128, 103, -23, -76, 127, -87, -27, 96, -55, -58, 60, 0, -95, 86, 49, -53, 42, -3, 45, -95, 54, 8, 1, -15, -48, -8, -55, 21, -39, 114, -90, 37, 91, -128, 91, -21, -18, -3, -13, -2, -55, 73, -128, 127, -90, -3, 58, -58, -8, -47, 29, -112, 87, -17, 33, 0, 0, 127, -100, 37, 36, -33, -58, 33, -1, -108, 119, -57, 7, -11, 23, -31, 60, -113, 66, 74, -118, 49, 54, -117, 127, -74, 24, -63, 107, -123, -2, 78, -128, 52, 8, -15, -65, 117, -128, 59, -16, 10, -22, 60, -6, 8, -65, 101, -39, -63, 111, -59, 50, -64, 106, -18, -60, 59, -121, 81, -75, 111, -116, 101, 24, -79, 95, -44, 43, -59, 65, -60, 34, 2, 21, 36, -10, 16, -10, 71, -112, 127, -91, 73, -85, 37, -70, 73, -65, -1, 88, -87, 45, -7, -44, 39, 22, -45, -17, 98, -128, 92, -75, -42, 93, -124, 57, 22, -86, 81, -78, 38, -58, 33, 38, -33, 90, -13, 45, -7, 86, -44, 98, -38, 31, -65, 65, -65, 12, -23, 13, 68, -107, -21, 127, -128, 127, -111, 48, 31, -92, 71, 37, -111, 78, 29, -58, 86, -10, 31, -10, 38, -34, -63, 92, -74, 52, -33, 57, 8, 70, -38, 65, 10, -78, 17, -13, -3, 36, -7, 57, 15, 63, -21, 48, 69, -76, -31, 36, -7, -111, 102, -2, -27, 64, -44, 63, -16, -10, 34, 3, 64, -74, 127, -49, -12, 1, 26, 34, -60, 123, -54, 6, 23, 53, -65, 95, 3, -64, 101, -102, 101, -128, 80, -2, -114, 127, -128, 63, -37, 81, -128, 127, -128, 106, -69, 68, -34, 75, -28, 55, -27, 87, -63, 23, -13, 49, -118, 93, -37, 3, -29, 68, -64, 85, -71, 63, 28, -100, 87, 6, -66, 75, 5, -49, -13, 37, -36, 3, -52, 79, 16, -100, 59, -63, 95, -87, 52, 34, -81, 31, -123, 92, -114, 96, -113, 127, -128, 108, -45, 0, 23, -16, 18, -96, 127, -106, 47, 36, -69, 1, 69, -39, 21, 23, 23, -47, -15, 52, -74, 22, 10, -16, 43, 12, -8, 8, -23, 24, -22, -36, 27, 69, -75, 91, 42, -78, 37, 60, -98, 70, -119, 127, -128, 122, -48, 0, -26, -59, 21, -47, -24, 28, -8, 17, -48, 47, -57, 54, -114, 78, -42, -66, 108, -42, -49, 52, -44, -17, 32, -90, 48, -8, -50, 86, -69, 15, 65, -128, 122, -66, -1, 87, -78, 97, -63, 1, 27, -91, 43, 60, -54, 73, -43, 26, 11, -10, -15, 85, 0, -6, -27, 27, -6, -60, 80, 8, -79, 118, -128, 127, -128, 109, -3, -53, 2, 87, -80, -7, 55, 10, 5, 8, 86, -102, 44, -24, -21, 13, -28, 93, -34, 52, -33, -52, 78, -128, 100, -3, -63, 107, -28, -28, 127, -128, 88, -55, 60, -127, 70, 0, -71, 91, -108, 93, -78, -36, 101, -79, -26, 63, -80, 58, -52, 58, -45, 18, -21, 11, -45, -78, 39, -32, -49, 33, 44, -49, 39, 15, -50, 18, 80, -55, 0, 100, -85, -65, 111, -113, -38, 63, -28, 7, 6, 33, -8, -22, 22, -39, -52, 127, -55, -22, 45, -42, 31, -54, 23, 55, -98, 2, 57, -109, 127, -128, 127, 0, -53, 55, -28, 66, -95, -38, 127, -128, 38, 34, -98, 91, -54, 10, 71, -78, 75, -37, 79, 0, -28, 122, -66, -28, 102, -122, 117, -128, 91, -3, -10, -16, 124, -128, 108, -12, -3, 37, 10, -54, 57, -91, -22, 13, 22, -101, 49, 27, 13, -78, 102, -43, 26, -74, -10, 13, 17, -44, 38, 5, 0, -68, 3, 81, -88, 117, -73, 37, 55, -128, 108, 7, -90, 91, 38, -128, 119, -71, -63, 107, -123, 54, -42, 50, -91, 127, -73, -43, 127, -103, -49, 127, -128, 108, -24, 8, -8, 27, 55, -7, -15, 73, 13, -75, 52, 12, -74, 38, 57, -98, 70, -74, 37, 0, -58, 96, -66, 31, 10, -39, 32, 8, 33, -49, 54, -50, 106, -128, 37, -10, 18, 13, -66, 28, 47, -128, 127, -96, 10, 27, -59, -21, -3, -23, -6, -3, -18, 32, 42, -128, 127, -22, 0, 34, -22, 80, -128, 45, 18, -93, 91, -23, -12, 73, -74, -15, 18, -75, 0, 10, 22, -69, 127, -57, -5, 42, -58, 27, -45, 26, -5, 12, 73, -45, -5, 5, 6, -79, 118, -121, 15, 106, -128, 118, -6, -88, 114, -128, 86, -36, 58, -55, 65, 63, -113, 81, -33, 6, 28, -38, 0, 114, -128, 101, -66, 3, 0, 53, -128, 127, -128, 127, -76, -11, 18, 5, -50, 11, -21, 106, -128, 33, 93, -128, 109, 18, -128, 127, -70, -28, 38, 27, -128, 127, -118, 65, -16, -27, 49, -53, -91, 81, -68, 12, -38, 65, 47, -100, 91, 49, -118, 111, -39, -21, 111, -90, 39, 28, -58, -22, -6, -63, 21, 18, 0, 53, -13, 38, -31, 79, -128, 124, -10, -60, 121, -17, -43, 107, -71, -33, 47, 29, -49, 73, 49, -95, 127, -128, 127, -74, -49, 88, -54, 76, -38, 63, -26, 54, -128, 58, -23, -33, 32, 58, -73, 88, 49, -119, 101, -34, 50, -45, 86, 11, -3, 32, 79, -108, 70, 1, -21, -26, 36, -75, -8, 44, -128, 127, -128, 127, -128, 75, -22, -17, 32, 26, -15, 79, -65, 44, -13, 39, 11, -96, 127, -128, 68, -10, -28, 38, -80, 45, 49, -118, 79, -3, 37, -59, 127, -54, -53, 81, -97, 47, -68, 122, -128, 86, 21, -31, 36, -11, 57, -74, -6, -12, 68, -128, 118, -113, 93, -80, 76, -107, 17, 49, -122, 107, -6, -6, -12, 24, 60, -128, 127, -85, -1, 101, -122, 107, 11, -96, 93, -12, -59, 13, 50, -119, 127, -128, 108, -49, 11, 37, -15, 23, 26, 1, -80, 127, -128, 127, -117, 6, 5, 7, -63, 87, -95, 103, -21, -96, 127, -80, 91, -78, 78, -33, -11, -13, 86, -128, 47, 0, -45, -23, 123, -111, -12, 127, -128, 65, 55, -97, 7, 0, 12, -102, 87, 22, -119, 96, 12, -103, 92, -57, 21, 6, -69, 71, -15, -6, 63, -57, 52, -24, 76, -111, 26, 39, -66, -1, -68, 85, -128, 92, -33, 13, -13, 37, 48, -15, 6, 32, -5, -45, 68, -53, 100, -15, 6, 26, -93, 127, -91, -49, 100, -98, 39, -55, 55, 37, -45, 34, -29, 92, -123, 52, -29, 60, -116, 70, -44, 29, 8, 11, 18, 18, -37, 34, -24, -53, 91, -59, -15, 2, 55, -69, 2, 57, -98, 118, -86, 63, -43, 17, 17, -16, -36, 53, 50, -59, 122, -1, -109, 124, -3, -100, 127, -91, 39, -13, 22, -68, 11, -49, 58, -47, -49, 127, -93, -3, -6, 33, -78, -50, 127, -91, -70, 127, -122, 12, 37, -36, 58, 6, 43, 10, -1, 5, -78, 52, -26, -18, 54, -38, 121, -128, 127, -97, 13, -21, 76, -114, 16, 27, -81, 31, -78, 22, -42, 28, 48, -92, 102, -34, -43, 37, -53, 93, -71, 34, -38, 65, -108, 15, 28, 37, -66, -3, 117, -128, 127, -96, 12, -10, 37, -128, 127, -128, 49, 5, -26, 1, 18, -24, 66, 22, -16, 53, 16, -97, 48, 8, -75, 17, 45, 8, -113, 118, -15, -5, 11, 85, -128, 116, -57, 0, -7, 87, -93, -3, 39, -39, 42, -21, -13, 116, -128, 13, 70, -91, 127, -107, 69, -6, -1, -27, -21, 76, -69, 18, -64, 47, -22, -78, 86, 64, -81, 47, 24, 12, -74, 47, -16, 7, -116, 91, -16, -128, 127, -128, -13, 78, -85, -5, 91, -98, 127, -113, 79, -43, -79, 116, -128, 34, 68, -128, 127, -44, -74, 127, -58, -47, 47, 12, -65, 11, 23, 5, -28, 48, -31, 3, 13, -52, -21, 59, -109, 43, -2, -21, -63, 37, -36, -37, 96, -128, 101, 31, -57, 26, 103, -123, 102, -96, 88, -55, 21, -58, 119, -119, 102, -71, 97, -128, 98, -52, 66, -34, -16, 127, -128, 127, -36, -64, 48, 11, -117, 93, 52, -109, 127, -100, 92, -44, -23, 15, 36, -128, 127, -63, -21, 54, 11, -37, 12, 18, -90, 88, -29, 44, -79, 93, -86, 31, -53, 78, 6, -78, 127, -128, 127, -113, 0, 39, -88, 42, -44, 88, -48, 10, 71, -128, 100, -13, -5, 17, 32, -78, 21, -59, 45, -50, 31, 50, -60, -64, 91, -76, -59, 92, 11, -68, 87, -7, -23, -66, 73, -127, 57, -69, 57, -57, -68, 127, -128, 54, -17, 45, -93, 114, -93, 88, -81, 42, -52, 85, -39, -28, 52, -24, -12, -29, 44, -60, 48, -39, -15, 68, -55, 66, -18, -11, 73, -128, 127, -128, 127, -39, -36, -3, 88, -128, 98, -36, 36, -69, 76, -102, 0, 26, -53, 55, -12, -71, 71, -27, -10, -37, 53, 8, -86, 101, -21, -86, 117, -114, 54, 0, 18, -15, 38, 18, -38, -27, 15, 66, -37, 15, 50, -21, -29, -10, 73, -106, 97, -128, 127, -101, 7, -54, 127, -128, 100, -65, 33, -22, 27, 29, -12, 43, 22, -1, -70, 127, -128, 22, 90, -128, 114, -52, 75, -85, 103, -3, -91, 127, -106, -24, 116, -112, 76, -32, -32, 12, -103, 38, -48, 12, 34, -2, 22, 5, 70, -57, 49, 71, -97, 39, -63, 32, 1, -116, 127, -122, 45, -31, 12, 11, -58, 127, -86, 8, 48, -27, -109, 100, -86, 76, -116, 127, -128, 112, -101, 57, 18, -106, 106, -63, 71, -36, 17, 103, -128, 127, -128, 78, 12, -60, 7, 116, -128, 119, -54, 1, 86, -95, 93, -12, -45, 70, -53, -28, 24, 11, -91, 117, -75, -24, 66, -74, 68, -128, 127, -28, -50, 116, -75, 88, 29, -21, 1, 50, -101, 32, -47, 24, -10, 42, -59, 64, -70, 8, 23, -10, 60, -16, 28, -47, 88, -43, 36, -55, 127, -128, 75, 22, -128, 127, -52, 5, 95, -80, 86, -34, -6, 7, -29, -15, 73, 2, -53, 32, 57, -102, 48, -3, -34, 81, -102, 53, 75, -128, 127, -118, 96, -127, 123, -80, 53, -48, 112, -100, 118, -128, 60, -16, 27, -55, 101, -39, 68, -66, 12, 6, -13, 23, -78, 92, 6, -53, 69, 18, -21, -10, 96, -69, -2, 68, -10, -80, 127, -106, 97, -69, 17, -23, 75, -88, 28, 48, -21, -79, 73, -57, -15, 81, -78, 76, -27, 33, -101, 49, -28, -13, -17, 31, -29, -15, -1, 33, -87, 64, -58, 18, -23, 97, -100, 79, -47, -3, -23, 53, 53, -80, 127, -102, 39, 0, -45, 58, -52, 13, -1, -3, -38, 45, 63, -78, 87, -15, 11, 0, -39, 13, -34, 5, 88, -111, 127, -101, 33, -31, 15, -79, 96, -87, 76, -7, -60, 53, -124, 117, -121, 2, 108, -128, 66, -12, -88, 60, -91, -29, 86, 5, -47, 103, -52, 52, -75, 32, 29, -76, -43, 69, -96, 10, 18, 79, -44, 33, 96, -92, -43, 127, -128, 114, -73, -15, 117, -128, 76, 11, -2, -16, 28, -6, -24, -11, 29, 1, -12, 49, -11, 24, -95, 78, 16, -2, -18, 59, -26, 49, -66, 59, 8, -16, 64, -2, -47, 31, -88, 76, -98, -1, 36, -86, 73, -128, 127, -128, 70, -17, -24, -33, -5, -63, 5, 34, 18, 32, 2, 8, -21, -33, 38, -64, 86, 33, -33, 18, 47, -36, -24, 76, -58, 3, 65, -86, -33, 85, -127, 95, -38, -24, 28, -90, 15, -5, 15, 1, -29, 87, -112, 12, -6, -24, -8, -17, 0, 49, -28, -31, 107, -55, -66, 127, -128, 43, 37, -37, -18, 127, -92, 11, 52, 0, -97, 97, -52, -75, 85, -71, 31, -60, 127, -78, 33, 59, -50, 108, -98, 127, -128, 70, -23, 5, 2, -6, 10, -42, 66, -128, 58, -21, 45, -78, 124, -92, 87, -73, 60, -31, 45, -80, 95, -85, 97);

    signal memory_control : std_logic := '0';      -- A signal to decide when the memory is accessed
                                                   -- by the testbench or by the project

    constant SCENARIO_ADDRESS : integer := 1234;    -- This value may arbitrarily change

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);

                o_done : out std_logic;

                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,

                o_done => tb_done,

                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;

    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.

        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;

    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_rst <= '1';

        -- Wait some time for the component to reset...
        wait for 50 ns;

        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench

        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock


        for i in 0 to 16 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_config(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);
        end loop;

        for i in 0 to SCENARIO_LENGTH-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+17+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);
        end loop;

        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component

        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));

        tb_start <= '1';

        while tb_done /= '1' loop
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;

        tb_start <= '0';

        wait;

    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;

        wait until rising_edge(tb_start);

        while tb_done /= '1' loop
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH-1 loop
            assert RAM(SCENARIO_ADDRESS+17+SCENARIO_LENGTH+i) = std_logic_vector(to_unsigned(scenario_output(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(17+SCENARIO_LENGTH+i) & " expected= " & integer'image(scenario_output(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(SCENARIO_ADDRESS+17+SCENARIO_LENGTH+i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done == 0 before start goes to zero" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;

