-- TB EXAMPLE PFRL 2024-2025

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity tb_gen4_mod5 is
end tb_gen4_mod5;

architecture project_tb_arch of tb_gen4_mod5 is

    constant CLOCK_PERIOD : time := 20 ns;

    -- Signals to be connected to the component
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);

    -- Signals for the memory
    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    -- Memory
    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

    -- Scenario
    type scenario_config_type is array (0 to 16) of integer;
    constant SCENARIO_LENGTH : integer := 5000;
    constant SCENARIO_LENGTH_STL : std_logic_vector(15 downto 0) := std_logic_vector(to_unsigned(SCENARIO_LENGTH, 16));
    type scenario_type is array (0 to SCENARIO_LENGTH-1) of integer;

    signal scenario_config : scenario_config_type := (to_integer(unsigned(SCENARIO_LENGTH_STL(15 downto 8))),   -- K1
                                                      to_integer(unsigned(SCENARIO_LENGTH_STL(7 downto 0))),    -- K2
                                                      1,                                                        -- S
                                                      11, -3, 5, 9, -4, 5, 10, -1, 5, -3, 2, 1, -3, 0   -- C1-C14
                                                      );
    signal scenario_input : scenario_type := (-104, 54, -17, 57, 93, -61, 112, -70, 9, -36, -11, -35, -114, 38, -22, -72, 61, 34, 121, -30, 108, 90, 62, -50, -111, -117, -50, -106, 43, -38, -48, -62, 105, -59, 58, -57, -49, -4, -50, -55, 9, -25, 65, -93, -17, -46, -111, -45, -74, 58, 61, 41, 5, 92, -98, -88, 61, 36, 113, 107, -4, 65, -3, 73, -85, -79, -120, -128, 37, -52, -111, 113, 122, 42, -23, 108, -47, 11, -29, -125, 88, 2, -68, -77, 93, 110, 10, -120, 117, 111, 55, -38, -10, 23, 4, 22, -95, 44, -27, -10, -121, -68, -88, -7, 92, 88, 80, -122, -46, 127, 36, -15, 46, -37, 51, 64, -38, 45, 62, -74, 40, 46, 30, 83, -57, -126, 104, -95, -71, -95, 48, 37, 35, 82, -7, 124, -62, -41, 81, 39, -78, 101, -49, -76, -71, -113, -74, -77, -106, 77, 58, -31, -116, 84, 65, 78, -33, -69, -121, -71, 58, 53, 77, -112, -32, -38, -7, 82, -11, -63, 33, 91, 65, 17, -48, 119, -16, -109, 45, 18, 24, -40, 123, -24, -32, -83, 99, -3, 76, -94, -108, -102, -2, -87, -46, 123, -33, 99, 27, -34, 81, -124, 32, 88, 16, -106, -10, -119, 32, -58, -54, 19, 87, -114, -115, 45, -7, -120, 37, 19, -5, 49, -76, 24, 117, -58, 5, -1, 68, -80, -4, 121, -37, 48, 63, 126, -65, 80, -89, 118, -58, 119, 125, 27, -105, -120, -103, -118, 96, 83, -106, 98, -3, -53, -28, -40, -91, 19, 22, -25, 25, -107, -128, 10, -6, -127, -49, -24, 19, -13, 118, -3, -82, 40, -70, -103, -81, 94, 48, -48, 71, 36, -15, 41, 7, 79, 104, 78, -104, -34, 54, -12, 87, -87, 82, 62, -51, -17, 30, -98, -111, -36, 2, 16, 103, -23, 56, 36, -11, 23, 127, -119, 56, -115, -65, 124, -5, -6, 17, 112, -71, -24, 39, 14, 54, 14, 123, 103, -13, -10, -47, -124, 38, 57, 22, 48, 47, -92, 3, 7, -16, -111, -28, 61, -49, -116, 76, -17, 112, -43, -115, 99, 34, 119, 40, 94, -22, -66, -35, -88, -70, 48, 57, 4, -11, 48, 8, -31, -83, 79, 21, -51, -123, -91, 114, 111, 123, 73, 96, 94, -124, 104, -35, -47, 28, 111, -44, 91, 22, -66, -103, -65, 80, -24, 86, 27, 4, -85, -11, -27, -1, 88, 44, -81, 105, 74, -67, -50, -20, 66, -63, -59, 97, 104, -18, 18, -13, -61, -30, -123, 30, -87, 79, 114, -81, -77, 18, -81, -23, 95, 58, 57, 91, 127, -3, -128, 63, -1, -94, 113, -39, 59, 69, 45, -68, 2, 126, 68, -50, 82, -63, 83, 39, -12, 69, 49, -60, -37, 119, -92, 94, -57, -26, -54, -65, -126, -91, 123, 35, -7, 4, 83, -37, 63, -74, 86, -120, -4, 10, 90, 65, 73, 39, -29, -77, -51, -91, -16, -127, 25, 104, 111, -126, -113, -44, -84, -35, 7, -98, 20, -71, -126, -77, -31, -91, -19, 39, 34, -116, 45, -93, -12, 28, -73, -56, 43, 34, 30, -54, -58, 116, -83, -77, -66, -7, 95, -111, -98, 125, -9, -6, -51, -94, -24, -13, 34, 28, -30, -106, -41, 76, -84, -115, 68, 94, 36, -2, -12, -39, -113, 115, 51, -9, 119, -47, -98, -40, 52, 105, 9, 70, 42, -4, 37, 88, 91, 40, -91, -96, -35, 114, 8, 56, 51, -55, -105, -106, -68, -73, 21, -126, -109, 127, 86, -26, 109, 124, -37, 50, -86, 19, -101, 79, -105, 15, 57, 110, 51, 108, 76, 2, -17, 47, 50, 12, -75, -69, 28, 86, 43, -3, -115, 10, -95, -48, 124, -101, 47, 65, -117, -105, -111, -110, 63, 15, -41, 79, 2, -65, 80, -12, 32, 88, -3, -49, -105, -54, -69, -97, -102, 111, -3, -41, 24, -102, -89, 52, -96, 72, 38, -88, -18, -101, 46, 90, 53, 33, 7, 59, -51, 7, 16, 4, -73, -81, -70, 125, 52, 45, 38, 118, 80, 18, -98, 119, -111, 30, -59, -111, 111, -113, 103, 11, -80, 126, 63, 81, 12, 103, -50, -2, 92, -32, 66, 24, 76, 101, 118, 79, 41, 59, -67, 120, 111, 60, 61, -66, -94, 48, 109, -81, 82, -110, -39, -15, 10, -58, 85, -28, -18, -102, -22, -105, 6, -18, 98, -47, 23, 124, -89, -14, -84, -47, -121, 109, -35, 87, -122, 42, 89, 115, 29, -112, 61, 113, 118, 119, 69, 114, 111, 70, -50, -74, 94, 42, 46, 114, 63, -128, 76, -18, -113, 12, -46, 115, 93, -47, 87, 57, 106, 108, -1, 100, -64, -60, -86, 78, -85, -123, 88, 31, 39, -69, 69, 52, -97, -73, 127, -33, 17, -75, 40, -44, 115, -127, 19, -2, 107, -57, -67, -96, -14, -4, 85, -75, 126, -77, 46, 35, 28, 109, 63, -106, -53, 90, 14, 25, -98, -40, -64, -29, -8, 100, 95, -87, -42, -44, 51, 18, -56, 94, -38, 97, -21, -62, -123, 18, -67, -55, 126, 30, 81, -16, 94, 107, -14, -92, -67, -58, 68, 42, -82, 64, 51, 53, 4, 88, 29, 89, -9, 17, -15, -72, 40, -40, 120, 43, -15, 92, -100, 114, -102, -61, 49, 126, 89, -79, 123, 56, 22, -16, 49, 87, -40, -1, -71, 113, 60, 46, -67, 38, -60, -4, -10, -90, -28, -47, -36, -12, 58, -85, 125, 43, 114, -39, -6, -81, 64, -119, 15, 106, -57, 119, 30, -39, -15, -89, -65, -70, -94, 103, 56, 35, -11, -68, 105, 69, -70, -126, 63, -61, 29, 90, 25, -17, 11, -90, 46, -62, -24, -83, 45, -35, 84, 86, 66, 97, 40, 61, 91, -56, 68, -43, 14, 42, 103, -38, 20, -8, 102, -125, 112, -9, 25, -90, 18, -91, 34, -73, -109, -86, -112, -105, 66, -109, -78, 81, 70, 86, 30, -84, 64, -7, -51, 18, 64, -116, 98, -53, -76, -77, 9, 85, 118, -47, 91, 68, -47, 126, -25, 0, 120, -10, 78, 126, -94, -50, 104, -54, 50, 115, 100, 41, 2, -117, -56, 115, -104, 9, 57, 79, -83, -126, 7, -25, 22, 71, -68, 14, -24, 95, 118, 126, -80, 18, 15, 32, 98, 27, -81, 35, 63, -99, -92, 71, 114, -67, -123, 69, 72, -83, -58, 57, 16, -5, -10, -72, 19, -76, -26, 97, 57, 115, -101, -126, 16, 4, -67, -101, -20, -51, -17, 100, 35, 18, 66, 72, -24, 47, -117, -40, -124, 77, 106, 15, -27, -26, 60, 78, -46, 28, 83, -107, 33, 101, 69, 26, 57, 126, -26, 32, 80, -94, 54, 107, -12, 82, 109, -74, 86, -36, 60, 93, 37, -25, -106, 113, -114, 69, 122, 11, 57, -101, -27, 52, 93, 13, -22, -15, -70, 120, 94, 104, -56, 118, 95, -56, 95, 62, -74, -107, 73, -64, 97, 24, -116, 86, -122, 32, 108, 98, 24, 99, 53, -114, 19, 37, -84, -60, -51, 91, 100, -120, 112, -16, 46, 40, 11, -63, 45, -63, 11, -30, 72, -19, -46, 31, -32, 111, -47, -109, -113, 35, -32, -60, 17, -14, -94, 122, 3, -32, -124, -67, 85, 42, -49, -96, 42, 27, -102, -23, 79, -20, 77, 81, -27, 1, 47, -49, -118, 7, -113, -70, -106, -100, 54, 69, -29, -51, 101, -60, -117, 21, 0, 39, -32, 26, 20, -42, 63, 76, 6, 122, -106, 13, -49, -80, -5, -72, -43, 121, 28, -90, -115, 46, 15, -39, 12, -58, -78, 69, -15, -34, -121, -24, -87, -109, 36, -36, 71, 72, -77, 109, -16, 79, -109, -91, -41, -13, 100, 67, 52, -46, -117, 110, -35, -19, 37, -72, -38, 17, -43, -12, -105, -116, -60, 7, 101, 71, -6, 20, 108, 22, 38, -71, 116, -94, 67, 113, -2, -121, 26, 44, 52, -89, -42, -98, 19, -40, 85, 6, 69, -104, -77, 52, -61, -11, -44, -86, 41, 26, 26, 105, -116, -104, 126, 17, -82, 75, 81, 107, 43, 100, 43, -56, 103, 39, -77, 46, -34, 7, -4, -99, 17, -115, 45, -112, 82, 47, -14, -82, 55, -118, 9, -68, 57, 73, 99, -18, 89, -87, -97, -95, -26, -48, 116, -27, 122, 48, 51, -47, 62, -42, 35, -23, 62, 2, -52, -82, 110, 115, 2, -16, 29, -128, 50, 60, -38, -20, 33, 68, -23, 126, -39, 22, 81, 120, 22, 79, -71, -4, -125, 105, -39, 105, 38, -39, 115, 6, -118, -47, -38, 25, -46, 111, -55, -109, 50, -84, -83, -32, -106, -53, -108, -119, -87, 38, 75, -56, -40, 108, -25, 16, 45, 35, 32, 119, -10, -103, -103, 84, -1, 56, 57, -69, -22, -62, 8, 121, -50, 53, -96, -91, -89, 92, -29, 124, -43, 104, -37, 67, 92, -104, -79, 26, 125, -81, 123, -70, 107, -20, 82, -38, 67, 96, 58, -34, -37, 123, 105, -115, 100, 66, 110, 51, -42, 97, -86, 119, 20, -1, 123, 100, 42, 18, 116, -122, 72, -57, 67, -16, 50, 103, -120, 32, 54, 89, -67, -81, 29, -128, -105, -107, -53, 102, 14, -100, -103, -72, -41, -106, 9, 15, -2, -57, 67, 48, 48, -92, 61, 91, -55, 11, 8, -124, -60, -16, -40, -16, 126, 71, 127, 108, 18, -20, -9, 27, 44, -93, 122, 100, 59, 121, -19, -12, -81, 82, -75, -127, 6, -45, -128, 77, 111, 95, 0, -31, 55, 31, -32, 89, 125, 62, -107, -36, -78, -127, -25, 119, -118, -113, -27, 50, 37, -27, 123, -53, -32, 63, 47, -122, 51, 73, -68, 82, -24, 47, 80, 2, -51, 57, 15, -39, 96, 55, -73, 11, -41, 70, -22, -37, 90, -94, 52, -32, 123, -21, -71, -58, -32, -54, 33, 99, -22, -53, 66, 86, 44, 71, 18, 71, 64, -25, 21, 45, -66, -30, -36, 43, -43, 99, -58, 10, 109, -71, -57, -14, 105, 127, -119, -53, 14, -27, -82, -108, -39, 105, 8, -69, 68, 118, 25, -118, -42, 1, 32, 87, -7, -98, -57, -85, 26, 61, 48, -26, 12, 113, 18, 40, 91, -92, -96, 43, -37, -62, 88, -59, 78, -22, -122, 115, -62, -44, 75, 11, -125, 35, -26, 65, -91, -27, -17, -37, -77, 93, -105, -75, 52, -119, 72, 39, -105, 32, 24, -63, -97, -37, -46, 78, 2, 62, -124, -18, 126, -49, 8, -12, -34, 113, -14, 43, 8, 93, -24, -47, -88, 5, -118, 3, 29, 57, 10, 22, 113, -101, 55, -109, 94, 117, -118, 15, -17, 32, 42, 120, -87, -110, 119, -12, 10, -103, -127, -3, 28, 81, 27, -95, -118, -50, -34, 103, -93, 87, -88, -60, 81, 36, -117, -44, 29, 33, -95, 101, -127, -116, 64, -24, 47, 111, -82, 105, 76, -115, -52, -81, 27, 9, -114, -77, -6, 16, 27, -99, 22, -82, -125, -12, 71, -9, -28, -76, -74, 47, -68, -44, 60, 13, 98, 33, 65, 97, -46, 5, 105, 111, -102, -60, 15, -106, -104, 26, 79, -123, 23, -44, -15, -22, -121, 49, -40, -103, -92, -59, -14, -61, -57, -24, 125, -59, 44, 108, 113, 119, -28, -75, 72, 78, 83, -14, 45, 84, 31, 109, 124, -50, -13, 99, -32, 102, 2, 125, -99, 110, -86, -22, 69, 103, 84, -3, 124, 120, -82, 6, 54, 44, 30, -5, -118, -54, -111, -77, -52, 25, 9, 87, 78, -15, 43, -18, 2, -28, 102, -33, 17, -39, 31, -53, 39, -90, -105, -54, -128, 86, 89, 13, -37, 123, 71, -104, 112, 88, -1, 97, -90, 87, 106, 120, -82, -21, 54, -6, -74, -102, -28, 105, 90, -27, 78, 2, 53, 105, 102, 8, 47, 97, -63, -65, 102, 24, 114, -13, -68, 38, -34, -57, 2, -118, -3, -33, 27, 23, 104, -98, -126, 80, -124, -60, 3, -80, -11, -124, -42, -117, -111, 94, 22, -100, -78, -77, -63, -58, -122, -121, -86, 32, 80, 107, -13, -38, 116, -5, 121, -9, 43, -17, 113, -37, -62, -103, 100, -115, 34, -47, 61, -42, 87, -61, 20, 22, -27, 41, 111, -119, -107, -63, -100, -4, 14, 52, 4, 125, -11, -44, 127, 94, 103, -37, -86, 2, 119, -14, -114, 96, 65, -76, -115, 33, 2, 27, 14, -27, 1, -77, 89, -22, -17, 43, 51, -2, -33, 58, -21, 16, 41, 24, 37, -46, -115, 124, 73, 28, 51, -91, 82, 91, 39, -7, -114, -84, 65, -83, 30, -13, -122, -93, -26, 27, -64, 51, -82, 4, -37, 53, -33, -49, -116, -73, 1, 34, -94, 61, 118, 68, 79, -72, 6, -26, -87, -64, 86, -89, 113, 92, -119, 110, 125, 74, -5, 41, -7, -117, 59, 54, 92, -9, -102, -125, -2, 73, 87, -76, 99, 71, -37, -60, 96, -55, -61, -46, 97, -76, 22, 29, -33, 15, -31, 75, -112, 104, 3, 61, 82, 127, 95, 39, -99, -8, -59, -17, 11, 81, -122, -43, -47, 124, 54, -22, -46, -24, 65, -78, 49, 28, -122, -70, -76, -46, 50, 45, 106, -19, 98, 40, -61, 28, 127, -34, -63, -29, 106, -61, -121, -123, 65, 11, -81, 75, -70, 66, -53, 127, -73, -100, 94, 62, 97, 127, 101, -4, 33, 82, 45, -37, 17, 116, 69, 120, -20, -21, -92, -60, -78, -22, 51, -90, 40, 70, -73, -72, 81, 31, -47, -37, -117, 52, 11, -13, 41, -12, -59, -50, 15, 55, 97, 49, 58, 74, -106, 43, 39, -45, -79, 10, 90, -84, -122, -120, -124, 96, 45, -17, -99, 81, -73, 40, 91, 33, -14, 32, 65, 124, 120, 67, 33, 80, -54, 55, -59, 99, 4, 114, -97, -9, -65, 85, 27, 60, -69, -8, 35, -54, -57, -113, 116, -118, -95, 87, 124, -46, -8, -62, -85, -55, 122, 126, 20, -119, -32, 63, -58, 11, -29, -87, 65, -85, -7, -108, 12, -115, 94, -36, 36, -64, -128, -88, 50, 80, -70, 103, -43, -80, -79, -11, -92, 96, 109, -45, 29, -87, 105, 85, 16, -107, -76, 93, -15, -38, 103, -55, -45, 124, -26, -44, 19, -84, -48, 23, -78, -22, -85, -15, 31, -63, -100, 72, -11, 40, -109, 90, 85, -124, 85, -69, 21, 58, -77, 75, 124, 113, 125, 110, -127, -43, -107, -107, 49, -69, -121, 40, 98, -119, 43, 25, -75, 6, -68, 78, 11, 44, -126, 53, -124, -54, -3, -2, -66, -19, 57, -21, -54, 75, -16, -59, -20, -16, 124, -64, 63, 108, 83, -39, -102, 0, -101, 35, -48, -19, 8, 88, 51, -45, 44, 40, -97, 45, 1, 71, -12, 6, 92, 9, 23, -74, 104, -60, 9, 76, -84, 33, -9, 103, -34, -113, -119, 28, 31, 94, -65, 87, -74, -70, 122, 8, 5, 0, 119, -23, 22, -69, -126, 95, -6, -85, 102, 111, -62, 2, -70, -5, 51, -88, 108, -67, -117, -16, -104, -16, 44, -51, 14, 66, -86, -4, 78, 100, 12, 43, 41, 123, -116, -16, -122, 71, 1, 56, -28, -92, -63, -12, 101, -14, -44, -108, -38, -114, 113, -116, -32, 15, 51, -49, 65, 63, -106, 11, -58, -66, -81, 56, -19, 14, 43, -110, 59, -108, -69, -62, -40, 5, 70, 96, 41, -101, -78, 111, 70, 99, -127, 60, 77, -41, 67, 24, 97, 124, -47, -39, -126, -83, 39, 41, -64, 95, 93, -120, 66, -61, -5, 113, 114, -13, -74, -121, -62, -17, 12, 81, -71, 8, 75, -78, -31, -21, 94, -8, 114, 113, 70, 1, 52, -104, -75, -12, 105, -52, 19, 66, -12, 84, 91, 58, 111, 8, 20, -57, 26, 8, 87, -118, 39, -118, 42, 107, 14, 30, -28, -56, 3, -64, 73, 96, 22, 72, -125, 46, 103, 93, 90, -71, -9, 82, 61, -46, -73, 88, 99, 117, 34, -104, 123, -67, 56, -116, 104, 123, 30, 20, -87, -28, -47, -49, 45, 11, -99, -110, 7, 64, -80, 82, 109, 40, 26, -103, -128, 14, -119, 63, 99, -115, 61, 36, -16, -5, -25, -22, -36, 17, -124, -46, -123, -40, 122, -20, 50, 36, -101, 52, 44, 81, 15, 75, -38, -113, -85, -27, 90, -63, 40, -51, -87, 74, -31, 46, -56, 16, 103, -123, -56, -45, -9, -91, 7, -56, 106, 10, -65, -125, -84, -42, 42, 81, 20, -30, 54, -89, -16, 33, -76, -72, 65, 119, 38, 96, 29, -4, 67, 89, 32, -36, 64, -22, -47, 103, -15, 47, -128, 81, 25, 30, -59, 127, -120, 85, -80, -111, 116, -97, 57, 27, 117, -23, 113, 26, -25, 66, 90, 80, 25, 105, 30, -122, 90, 52, 32, 90, -27, -10, 88, -24, 92, -68, -27, 8, 57, 28, 72, -106, 110, -54, 109, 35, 127, 19, -81, -73, 3, 99, 31, 81, 92, -49, -4, 70, 55, -1, 10, 44, 80, 97, 106, 77, -53, -12, -28, 45, 73, -28, 119, 62, -93, -84, 97, -113, 63, 83, -123, -23, 81, -3, 125, 100, 13, -20, 97, 51, 15, 36, -7, 35, -102, 110, 22, 13, -39, -85, -64, -108, -56, -82, -81, 86, -12, -81, 14, 87, -106, -83, 75, 103, 111, 21, -116, 123, -128, 67, 81, -47, 19, 110, -115, -21, -13, 92, 70, 72, -128, -101, -95, 29, 44, 44, 122, -91, -91, -48, -15, -41, -43, -114, -73, 38, -25, -58, 106, 84, -57, -21, -92, 64, -56, 2, -53, -97, 47, 79, 11, 62, 127, -27, -79, -2, 110, -58, 4, 127, 105, 0, -45, 124, 50, 82, -65, 97, 7, -42, -106, 92, 64, -34, 15, -128, 34, -23, -97, -42, 93, 79, -12, 92, -44, -106, 48, -109, 91, -53, 46, 98, -52, 31, 10, 37, -69, -5, 37, -100, -104, 101, 17, -9, -95, 86, 112, 94, 49, -55, 70, 35, -80, -92, -10, -70, -11, 7, 123, 8, -77, -103, -24, 95, 66, -6, -113, 19, -81, 52, 44, -74, 35, -83, -97, -120, -57, -105, 34, -26, -93, -110, -71, 12, -112, 112, -58, -83, -12, 122, 126, -25, -80, -7, 72, -87, 61, -114, 68, 27, 61, -79, -70, -83, -69, -61, -62, 121, 84, -128, 31, -66, -26, 96, 47, -17, -8, -99, -128, 29, 0, 6, 45, 74, 126, 30, 31, -123, -18, -22, 86, 44, -4, -42, -67, -71, -32, -128, -76, 78, -20, -104, 75, -107, 59, 28, -37, -111, -87, -43, -95, -91, 60, 74, -36, 81, -5, 105, -26, -44, 83, -103, -16, 32, -109, 125, 59, 73, 49, -128, -45, -12, 8, 0, 73, -118, 115, -21, -49, -105, 127, -104, -62, -50, -69, -67, -1, -33, -68, -42, 76, 40, 122, -66, 113, -72, -16, -43, -96, 58, -13, 19, 74, 21, 84, -26, -95, -96, -128, -4, -75, 97, 120, 37, 103, -123, 91, -2, -66, 51, 85, 53, -16, -13, 52, -127, 89, 87, -108, -42, 91, 70, 49, -94, -95, 7, -94, -104, 80, -123, 2, 3, -89, 44, 87, -23, -122, -106, -37, -29, 87, -54, -96, 33, 15, 51, -21, 108, 17, -49, -111, 26, -36, 17, 74, 73, -81, 86, 27, -95, -19, 60, -73, 20, -66, -66, -12, -24, 96, -118, -87, 76, -61, 86, 25, 2, -72, 82, -103, -106, -44, -89, 6, -101, 24, 17, 23, 22, -128, -44, 33, -68, -108, 120, 124, 121, 11, -94, 65, 120, 26, 72, -103, 5, -76, -126, 93, -86, 87, 25, 46, 123, -101, 75, -27, -128, 77, -103, 38, 25, 27, -94, -89, 64, 127, 2, 108, 103, -87, -119, 118, -37, -62, 120, 117, -85, 40, -9, -101, 47, -35, -18, -48, 95, -43, 117, -76, -102, 36, -108, 110, 42, 113, 23, 123, 56, 121, -45, 65, -47, 97, 13, -62, -54, 79, 124, -97, 84, -90, 38, 51, -115, -41, -85, -43, 86, 38, 56, -86, -70, 15, 97, -105, 65, 34, 22, 70, 1, 39, 89, 88, -94, 18, 97, 3, -12, -105, -3, 34, -19, -43, 25, -50, 96, 112, -43, 104, -71, 29, -98, -79, 51, 88, 7, 120, -64, 66, 19, 115, 76, 44, -44, 126, 14, 25, 60, 91, -31, -37, -48, -64, 62, -72, 117, 69, -31, -57, 6, 59, -83, -5, -61, -126, 20, 0, -62, -50, 65, -79, 52, -121, -6, -29, -104, -34, 44, -73, -6, 67, 103, 92, -4, 33, 7, 123, 2, -14, -37, 20, 2, -70, -91, -24, -85, 121, -30, 96, 100, 102, 112, 38, 85, 123, 93, 4, -69, -15, 88, -127, -128, -104, -79, -62, 73, -30, 5, -46, -119, -84, 55, 51, 33, 25, -103, 37, 16, -3, 85, -17, 99, -89, 112, -67, 45, -59, -109, -96, 47, -8, 17, 123, 58, 127, 61, -46, -61, -9, -12, 18, 95, 29, 59, -90, 118, 0, -15, -41, 121, -88, -55, -87, -11, -31, -41, 79, -126, -84, -106, 35, 13, 102, -32, 99, -54, 79, -64, 93, 4, 95, -45, 52, 27, -99, 52, 100, -41, -94, -90, -98, -124, -123, 86, 3, 83, 8, -18, -41, -69, -50, 15, -58, -96, -1, 87, -72, 17, -13, 24, 67, 114, -107, 7, 48, 29, 67, 118, -102, 19, -15, 70, 60, -23, 63, -89, -27, 77, 78, 24, 32, -97, 98, 97, -46, 44, -96, 17, 74, 100, -87, 12, 6, 118, -47, 84, -68, -52, -12, -110, -9, 116, 12, -4, 44, 96, -36, 116, -70, -127, -121, 67, -8, -98, 10, -76, 105, 122, 68, -77, -101, 115, 24, 48, 81, 81, -2, -6, -11, -28, -54, -40, 37, 20, -31, -90, 12, -10, 52, -2, 104, -80, -104, -115, 59, -7, 115, -16, 78, -2, 3, 110, 40, -52, -50, 98, -8, 3, -7, 97, 3, 50, 21, 15, 100, 80, -109, -119, 54, 112, 93, 0, -6, 84, 122, 77, 28, 116, -65, -22, 21, 11, 35, 21, 42, 64, 88, 108, -70, 105, -118, -61, 53, 67, -54, -26, -62, 75, -38, 58, 101, -87, 60, 27, -4, 64, -59, 11, -46, -101, 39, -45, 33, -70, -88, 21, -124, 123, -48, -57, -28, 43, -117, -70, 5, -5, 39, -17, -41, -16, -87, 61, -17, 8, -79, 114, 56, -64, -85, 78, 45, -6, 4, -30, -108, 44, 80, 18, -34, -33, -91, -90, -49, -64, 28, -94, -97, -31, 119, 17, 103, -37, 39, -26, 81, -57, -77, -63, 42, 0, 11, 17, 63, -81, 107, -26, -31, 10, 117, -15, -94, 114, 88, 37, 46, 74, 2, 37, 10, 119, 86, -73, -80, -59, -119, 10, 14, 124, 46, -107, -71, -23, 15, 9, -49, -16, 17, -123, -42, 36, 124, 114, -45, -115, -16, 54, -17, 29, -8, 56, 39, -62, -31, -26, 108, 103, -109, -117, -73, -115, 66, -46, 117, 113, 113, -53, -114, 81, -43, -88, 39, -128, 25, 44, 89, 57, 72, 109, -51, 58, 8, 60, 97, 8, -120, -34, 31, -51, 20, -26, 126, -10, 58, -4, -86, 15, 45, -87, 88, 25, -64, -111, -92, -23, 127, 94, 2, -68, 94, -41, -6, -18, -4, -65, 71, -44, 19, 100, -59, 95, 41, -56, -37, 104, 65, -56, -74, -121, -49, 40, -18, 125, 109, 20, 91, 97, -49, -50, 18, -88, -43, 26, 87, 64, -76, 127, -61, -3, -95, 81, -10, 62, 74, 13, 9, 49, 115, -40, 94, -83, 79, -8, 77, 54, 31, -102, 58, -98, -20, -98, -84, 79, -95, -18, 93, 102, 52, -58, 118, 45, -119, -62, -55, 53, -14, -102, -42, 39, 43, -68, -29, 53, -24, -84, -94, -36, 19, 4, 127, -19, 80, 109, -44, -1, 77, -96, -110, 59, -4, -20, -15, 52, 23, 106, -115, -36, -116, 59, 37, -118, -128, -93, 105, -114, -38, -77, 59, -86, -59, -106, 60, -112, -30, -80, -103, 53, 25, -82, 41, -111, -72, -3, -60, 85, -25, -35, 75, 4, 59, 43, -25, 6, -115, 51, 27, -106, -92, 101, -69, -13, -121, -49, 63, 45, -9, -29, 57, 81, -124, -71, 37, 120, 27, 24, -24, -60, -84, -85, 33, 13, -90, -75, 77, -62, 32, 94, -52, -71, -53, 46, 3, -92, 85, -105, -49, -33, -33, 28, -6, 53, 93, -108, 105, 95, 16, 105, -119, -106, 116, -67, -72, 46, 76, -85, 37, -120, -29, -20, -21, -36, -128, 55, -82, 65, -114, 105, -103, 32, 99, -6, -127, 10, 95, 33, -16, -24, -82, -5, 110, 103, -74, -25, 104, 99, -47, -84, -101, 71, -124, 54, 45, -26, 27, 32, 99, -106, 87, -93, 58, -12, 39, -22, -62, -80, -70, -68, 83, 112, -123, 120, 23, -11, -100, 46, -39, 6, 25, -90, 119, -15, -48, -47, -48, 113, -47, 7, 75, -53, -120, 76, -29, 107, -110, -12, -110, -34, 108, 31, -111, -69, 122, -99, -93, -117, -121, 113, -19, 74, -34, -101, 112, -44, -85, -120, 90, 95, 7, 27, 87, 55, 80, -101, 5, -99, -6, 53, -76, 81, -43, -99, 3, -90, -3, 110, 4, -41, 78, -55, -61, 122, 94, 54, 15, 73, 79, -63, 108, -94, 12, -72, 112, 100, -125, -20, 51, 121, 61, -60, -55, 6, -48, 88, 91, 9, -1, -120, 63, -48, -119, 116, -81, 58, 29, -90, 121, -90, 35, 67, -103, -103, -29, -88, -58, 24, -74, 88, 122, -39, 8, -109, 95, -43, -120, 1, -59, 68, 70, 51, 33, -48, 87, -4, 26, 106, -42, -38, 27, -11, -62, -113, -117, -80, -80, -58, -78, -92, -113, -119, -9, 45, -55, -58, 34, 100, -80, 87, -9, 125, 40, 72, 31, 26, -2, 26, 113, 58, 26, -122, -56, -28, 50, 74, 25, -19, -127, -56, 125, 45, 98, 8, 15, 122, -55, 101, -83, -117, -116, 63, -6, -80, -45, -35, 88, -42, 23, -14, 116, 79, -124, 24, -53, -83, 74, -54, -100, -85, -11, -59, 69, -29, 20, 2, 49, -53, -6, -123, -90, 98, 93, 115, 27, 81, 61, 8, -111, -96, -79, 11, 51, 43, 12, 115, 113, 8, -109, 16, 67, 44, -109, -5, 89, 92, -70, 38, 39, 50, 119, -25, 122, -56, 29, -110, 40, -98, 78, 110, 73, -79, -52, -8, 69, -15, -95, -38, -72, -63, 36, -70, -70, 97, 12, 58, -27, 99, 124, 40, -37, 126, 92, -92, -128, 8, 69, -113, 116, -30, 32, 85, -96, 8, -36, -30, 102, 75, -63, 103, 64, -98, 61, 16, -35, -50, -6, 125, -63, -65, 54, 42, 120, -97, 27, -117, 54, 98, -39, -37, 32, -11, -92, -12, 14, -125, -42, 97, 27, -89, -9, 18, -34, 50, 103, 15, 44, -46, -34, 34, -5, 116, 68, 78, -24, 21, -115, 94, 28, 90, 104, -12, -4, -29, -114, 84, -93, -35, -30, -128, 23, 84, -62, 29, 67, 93, -98, -65, -33, 8, -28, 6, -37, -25, 25, -119, -45, 57, -126, -68, -79, 108, -9, -20, 8, 58, -121, -28, 105, -95, 74, 50, 31, -97, 66, -94, 67, 63, -118, 116, -110, 33, -111, 2, -112, 89, 53, 48, 119, 113, -53, -74, -24, -68, 90, 10, 101, -46, 103, -44, 15, 15, -17, 26, 81, 64, 90, 125, 17, 126, -121, -52, -52, -51, 15, -113, 98, 99, 63, -123, 9, 22, 68, -85, -85, 65, -91, 43, 84, 39, 58, 2, 23, -17, -100, -104, 69, -80, 16, 96, 118, -51, 22, -95, 58, -79, -30, -18, 53, -11, 44, 4, 110, 123, 119, 100, -126, 61, 115, 125, 33, -34, 27, 114, -85, -106, -111, -115, 65, -92, 73, -38, 85, -90, -127, 117, 34, 93, 74, -15, -77, -32, 102, 22, -127, 96, 49, 13, -105, 79, 61, 6, -93, -29, 51, 68, 35, 57, -117, 48, -67, 58, -23, -123, -47, 101, -16, 74, 80, 17, 18, 3, -58, 62, -13, -33, 127, 66, -36, 19, 6, 61, 101, 0, 110, -57, 103, -54, 120, -78, -99, 83, 73, -119, 81, -62, -3, 109, -3, -29, 127, -114, -17, -7, -27, -14, -67, 93, 117, -120, -93, 30, -48, 70, 122, 33, -57, -97, -58, 81, -59, -80, -63, 7, -128, 121, -52, -59, 36, -20, -101, -24, 71, -101, 94, -84, -20, 21, -79, 4, -28, -41, 22, -49, 100, -89, 119, -101, -104, 62, 126, 93, -52, 99, 15, -79, 101, 120, -91, -54, 107, -7, -126, -34, 50, -42, -114, -67, 121, -39, -13, -51, -108, 109, 82, 3, 48, 31, -116, -18, -33, 86, -66, -54, 61, -67, -81, 60, 30, -2, -77, 45, -15, 42, -14, 39, -119, 62, 22, -114, 79, 30, -40, 90, 3, -54, -97, -78, 47, -112, 51, -106, 21, 97, 26, 127, 6, -9, 119, 115, 62, -76, -12, -13, -16, 118, 19, -110, -7, 83, 33, -11, 112, -87, 118, -100, -115, -84, 70, 56, 91, -25, 14, 22, -85, 54, -62, 29, 83, 21, -62, 126, 38, -46, -49, -67, -22, 122, 96, -57, -124, -42, 47, -102, 58, 76, -116, -40, -28, 6, -59, 87, -36, 115, 99, -56, -27, 22, 39, -76, 118, -90, -98, -5, -86, 72, 83, -96, -114, -122, -126, 50, -17, -97, -69, -27, 67, 36, -117, 33, 51, -89, 9, -125, 9, 79, 37, 30, 74, -110, 43, -73, 123, 19, 21, -57, -31, 78, -73, 34, 63, -89, 114, -27, 118, 74, 15, -16, 0, 121, 88, -95, -66, 30, -120, -92, 49, 27, 42, -97, -61, 65, 61, 85, -117, -84, 127, 66, -94, -75, 32, 11, -90, 117, 91, 36, 127, 99, -55, -123, 7, -119, 126, -72, -26, -49, 55, -12, -98, -21, -86, 84, 29, -19, -112, -127, 90, -126, -47, 52, 86, -2, 32, -31, -14, 62, -107, -57, -74, 92, -87, -48, -80, 9, 113, 69, -35, 85, -84, 69, 38, 68, -23, 25, 70, -25, -80, 77, -117, 28, 19, -46, -41, 121, -119, 92, -66, 46, 28, -56, 60, 127, -24, -43, 34, 113, -41, -108, -34, 76, -35, -53, -74, 59, -42, 72, 66, 113, 19, 101, 98, 106, -118, -92, 58, 46, -81, 65, -70, -127, -112, 84, 13, -11, -97, 85, -72, -79, 22, -84, 81);

    signal scenario_output : scenario_type :=(-1, 3, -14, 12, -8, 3, 11, -11, 13, -7, 7, -7, 0, 7, -14, 2, -2, -3, 2, -7, 12, -3, 11, 4, 2, 0, -7, -5, 5, -8, 0, 1, 0, -7, 15, -11, 8, -1, -5, 2, -4, 0, 4, -6, 13, -8, 1, -3, -10, 2, -5, 0, 8, 7, -11, 8, -7, -10, 9, -3, 4, 5, 0, 9, -2, 11, -11, 0, 3, -19, 0, 4, -7, 0, 8, 4, -7, 17, -12, 0, 9, -10, 1, -4, 2, 0, -3, 0, 7, -8, 7, 1, 4, -3, 3, -1, -2, 7, -5, 7, -3, 2, -13, -2, -4, 6, 5, -8, 9, -3, -8, 10, 0, -7, 9, -6, -1, 11, -7, -2, 8, -10, 7, 9, -10, 10, 5, -13, 8, -9, 0, -10, 6, -2, 2, 11, -14, 10, 1, -10, 6, 11, -10, 13, -2, -2, 2, -11, -5, 4, -3, -1, 0, 2, -7, 10, 3, 5, -8, -2, -6, 1, 5, -2, 9, -13, 2, 3, -6, 1, 0, -3, 3, -2, 3, 11, -13, 7, 2, -7, -1, 1, 8, -6, 4, -3, 1, -5, 15, -5, 5, -2, -1, -15, 7, -5, -8, 17, -12, 13, 1, -14, 14, -4, 0, 7, 1, -8, 9, -14, 1, 4, 2, -9, 9, 2, -13, 1, 6, -12, 8, 0, -10, 12, -5, -4, 8, -1, 2, -11, 12, -6, -8, 7, 0, 0, 1, 7, -9, 8, -20, 18, -2, 9, 6, 5, -12, -8, 8, -15, 3, 15, -13, 9, 3, -6, -3, 3, -8, 6, 7, -9, 3, 3, -8, 0, 2, -7, -5, 0, 9, -10, 10, 6, -8, -1, -4, 2, -11, 4, 8, -8, 4, 0, -7, 3, 5, 3, -3, 9, -10, 1, 2, -10, 17, -10, 1, 10, 0, -5, 3, -4, -9, 2, 0, -5, 11, -6, -2, 10, -3, -1, 19, -25, 11, -2, -10, 5, 3, 2, -8, 11, -7, -1, -1, -4, 9, -2, 6, 11, -7, -4, 3, -10, 1, 9, -1, -1, 8, -2, 0, -5, 6, 0, -10, 5, -2, -8, 17, -15, 7, -1, -11, 7, 0, 12, -3, 9, 0, -9, -1, 0, -3, 0, 3, 3, 0, -2, -1, 6, -4, 7, -7, -4, -5, -8, 5, 0, 14, -4, 1, 17, -20, 5, 2, -5, -3, 17, -4, 6, -4, 0, -5, -7, 11, -2, 5, 0, 3, -11, 1, 5, -8, 0, 13, -8, 4, 2, 0, 1, -11, 3, 2, -6, 3, 10, -3, 5, -2, -2, 0, -18, 17, -5, -2, 13, -4, -12, 4, -4, -6, 2, 5, 9, -4, 5, 10, -20, 7, 3, -17, 12, -1, 2, -5, 4, 1, -7, 9, 3, -11, 13, -12, 4, 8, -2, -4, 10, -5, -6, 18, -13, 12, -1, 1, -11, 0, 0, -10, 5, 4, -2, 0, 4, -2, 9, -15, 9, -11, 1, -2, 8, 4, 3, 4, -1, 0, -2, -14, 3, 0, 5, -1, 12, -7, -8, 5, -6, -1, 11, -9, 2, 1, -6, -7, 1, 1, -4, 3, 8, -17, 13, -5, -5, 3, -3, -1, 5, -7, 8, 3, -9, 10, -11, 4, 2, -14, 12, -1, -9, 15, -4, 0, -2, -6, 3, 3, 0, -4, 6, 0, -12, 3, 0, -7, 4, 6, 5, -8, -3, 7, -18, 12, 10, -8, 5, -6, -2, -3, 0, 10, -4, 0, 0, 0, 6, 6, 1, -2, -2, -3, -7, 14, 1, 3, 3, -1, -6, 0, 3, -18, 3, 1, -15, 2, 13, -7, 6, 9, -4, 3, -5, 7, -18, 8, -9, 0, -1, 9, 0, 1, 2, 1, 1, 4, -2, -2, -2, -2, 5, 1, 3, 5, -19, 12, -5, -13, 24, -6, 2, 9, -13, -4, 2, -13, 5, 7, -11, 6, 2, -12, 10, 1, 2, 5, 0, 2, -3, -9, -1, 3, -13, 14, 3, -11, 9, -7, -11, 17, -11, 7, 1, -13, 5, -7, 2, 2, 4, 2, -4, 7, -1, 3, 0, -5, -4, 0, -9, 4, 0, 5, 4, -1, 7, 5, -13, 22, -21, 10, -2, -15, 23, -23, 5, 4, -9, 6, 3, 7, -11, 13, -6, -4, 7, -9, 2, -1, 3, 1, 9, -2, -6, 9, -10, 11, 9, -5, 0, 5, -10, 4, 14, -15, 10, -5, -5, 0, 6, -5, 7, -1, 1, -8, 0, -4, 4, -13, 17, -3, -2, 13, -5, -4, -4, 2, -7, 10, -15, 10, -9, 10, -2, -1, 3, -12, 3, 1, 0, 6, 5, 7, -3, 3, 0, -12, 6, 10, -5, 3, 17, -18, 7, -3, -13, 12, -11, 2, 6, -10, 9, -3, 6, 11, -5, 3, -1, 7, -19, 7, 0, -7, 4, -4, 13, -5, -6, 8, -2, -7, 10, -5, 0, -1, 7, -13, 11, -8, 9, -3, 8, -6, -4, -1, -3, 0, 10, -17, 15, -13, 2, 10, 0, -3, 7, -4, -1, 8, -2, 5, -8, -4, -6, 7, -1, 2, 5, -7, 4, -9, 5, 1, -7, 15, -4, 4, 0, 3, -19, 5, -2, -6, 7, -7, 11, 0, 3, 6, -4, -6, 5, -9, 0, 6, -7, 1, 0, 2, -1, 7, -2, 10, -6, 2, -3, -8, 11, -12, 13, -1, -2, 17, -22, 8, -7, 3, -5, 1, 12, -10, 6, -2, 6, -1, 2, 1, -7, 6, -5, 5, 2, 6, -9, 10, -5, 0, 3, -7, -2, 2, -6, -5, 7, -8, 12, -1, 5, 0, 3, -18, 17, -14, -3, 17, -10, 11, 3, -3, 4, -12, -4, 2, -8, 11, -5, -1, 9, -3, -1, 6, 0, -18, 10, -3, 0, 9, -1, -1, 6, -7, 3, -4, 0, -12, 7, -8, 4, 3, -2, 10, -2, 1, 9, -12, 4, 0, 1, -2, 4, 1, -1, -7, 17, -12, 9, -1, 3, -7, 12, -8, 8, 0, -11, 3, 1, -18, 7, -6, -6, 11, -3, 2, 9, -11, 2, 7, -9, 0, 15, -13, 7, -8, -5, 1, -3, -2, 17, -14, 6, 9, -18, 14, -3, -10, 19, -1, -8, 15, -6, -13, 10, -4, 3, 10, 4, -8, 9, -4, -13, 12, -3, 6, -4, 6, -3, -12, 8, -2, -1, 4, -11, 2, 2, 4, -1, 11, -12, 3, 6, -4, 0, 11, -3, -6, 1, 2, 0, -5, 4, 5, -8, -2, 6, -2, -5, 7, -1, 1, 3, -13, 4, -6, 2, 13, -8, 8, 0, -5, 0, 2, -1, -12, 1, 0, -6, 4, 4, -2, 6, 7, -3, 2, -15, 7, -7, 4, 2, -2, 4, -4, -3, 14, -6, -8, 10, -8, 0, 0, 7, 0, -5, 17, -6, -7, 14, -11, -3, 15, -8, 2, 10, -17, 11, -2, 6, -3, 6, 0, -22, 20, -12, 7, 9, -9, 4, -5, 1, 0, 8, -6, -5, 2, -3, 2, -3, 18, -13, 2, 15, -4, -2, 7, -4, -12, 20, -15, 10, 5, -22, 12, -8, -1, 3, 14, -5, 0, 13, -7, 0, 0, -9, 9, -11, 1, 13, -18, 12, 0, 0, 3, 3, -7, 3, -5, 7, -8, 7, -5, -1, 12, -6, 4, -1, 0, -11, 5, 4, -12, 1, 8, -7, 11, -9, 0, 0, -2, 0, 0, 6, -8, -3, 7, -8, -7, 12, -4, 0, 9, 2, -5, 7, 2, -8, 8, -13, -4, 1, -4, -3, 8, 6, -12, 8, -1, -7, 2, -3, 7, -7, -2, 6, -9, 9, 6, -7, 18, -13, 5, 0, -13, 3, 4, -3, 2, 0, 1, -10, 6, 5, -10, 3, 2, -3, 5, 0, 6, -13, 2, -4, -12, 13, -10, 2, 7, -6, 15, -9, 8, -11, -5, 0, 0, 11, -7, 4, 4, -17, 15, -1, -6, 7, -3, 0, 7, -5, 0, -9, -6, 1, -2, 0, 5, 0, 1, 1, 2, 4, -19, 19, -3, -1, 2, 2, -4, 4, 1, 3, -6, -1, -8, 4, -1, 11, -10, 11, -4, -6, 11, -9, -1, 1, -11, 11, 6, -14, 11, 2, -17, 5, 1, -7, 2, 1, 11, -7, 3, 11, -12, 7, 5, -9, 11, -6, 3, 0, -6, 4, -15, 14, -8, 1, 6, 1, -9, 7, -15, 4, -3, 0, 5, 13, -6, 8, -4, -8, -3, 0, -9, 13, -5, 5, 0, 5, -7, 5, -5, 8, -2, -2, -4, 4, -6, 2, 13, -4, -8, 12, -10, 0, 2, 0, -6, 2, 8, -13, 8, -2, -1, 5, 8, 0, 2, -7, 4, -15, 18, -14, 7, 12, -8, 6, 0, -5, -5, 0, 12, -14, 13, 3, -12, 11, -3, -2, 6, -6, -4, -7, 1, -3, -6, 9, -1, -9, 9, -3, -4, 4, 8, 0, 0, 0, -3, -12, 14, -2, 2, 4, -12, 6, -4, 0, 17, -8, 0, -4, -4, -6, 8, -7, 11, -14, 19, -2, -4, 3, 0, -8, 0, 10, -13, 13, -9, 9, -11, 9, -1, 4, -3, 0, 9, -11, 0, 10, -13, 12, -5, 9, 0, -10, 17, -19, 6, 3, -3, 1, 12, 0, -4, 12, -14, 9, -13, 15, -4, -6, 10, -6, 7, -5, 13, 1, -7, 7, -14, -1, 3, -3, 6, 1, -1, -6, -5, 3, -4, -2, -1, 2, 0, 1, -5, 13, -9, 0, 15, -5, -2, 6, -7, -9, 0, -3, -7, 11, 2, 4, 3, -1, 4, -7, -5, 9, -15, 10, 7, 0, 3, 0, 10, -14, 9, 4, -17, -3, 2, -7, 7, 0, 4, 3, -8, -2, 4, 2, 3, 5, 11, -10, -7, 7, 0, -9, 8, -7, -2, -7, 6, 7, -13, 10, 3, -7, -3, 14, -15, 2, 8, -14, 11, 0, -3, 4, 5, -11, 2, 9, -7, 5, 2, -6, 7, -12, 11, -2, -7, 7, -9, 13, -8, 9, 0, -5, -7, 4, 0, -5, 3, 0, -6, 3, 2, -2, 8, -2, 0, 9, -2, 0, 2, -2, -3, -1, 7, -15, 17, -1, -5, 4, -9, 8, 0, -2, 13, -4, 0, 0, -7, 0, 1, -10, 1, 5, 0, 1, 2, 2, -11, 1, 6, 0, 6, -1, -9, 0, -3, 1, -3, 5, -1, -7, 14, 3, -7, 10, 0, -14, 8, -2, -7, 19, -18, 8, 7, -21, 13, 3, -9, 3, 3, -7, 7, -8, 10, -4, -6, 4, 5, -17, 18, -9, -11, 19, -15, 1, 11, -5, 1, 2, -6, -5, 0, 0, 7, -14, 14, -7, -6, 14, -12, 3, 1, -7, 7, -2, 7, -1, 5, 1, 0, -11, 5, -8, 1, -5, 10, -1, 0, 8, -20, 22, -12, 0, 11, -13, 0, 4, 8, -12, 11, 0, -8, 17, -8, 0, -5, -7, 7, 3, 2, 2, -9, 0, -2, -4, 18, -21, 10, 3, -5, 0, 4, -1, -8, 5, 13, -22, 13, -6, -15, 14, -7, -5, 22, -10, 5, 5, -10, 7, -4, -1, 2, -6, 1, -1, 1, 11, -13, 0, 0, -4, 0, 7, -6, 3, 0, -12, 6, -6, -4, 5, -7, 11, 0, -6, 5, 4, 0, -1, 15, -3, -9, 0, 4, -8, -1, 12, -12, 10, -7, 0, 9, -9, 5, -2, -2, -1, -4, -5, 2, -1, -13, 10, -9, 6, 9, -3, 3, 0, -4, 3, -2, 7, -6, -3, 12, 0, -4, 12, -7, -4, 6, -2, 5, -4, 18, -22, 9, -7, 1, -2, 0, 14, -5, 0, 10, -7, 1, 8, 1, 2, 4, -8, -1, -5, -4, -6, 6, -3, 4, 6, -3, 0, 0, 3, -5, 8, -3, 1, -1, 10, -8, 9, -10, -11, 6, -8, -1, 2, 11, -13, 1, 13, -17, 11, 2, -12, 10, -3, 6, -4, 12, -2, 0, 2, -6, -4, 0, -6, 4, 6, -11, 4, 0, 0, 0, 11, 1, -8, 8, -5, -5, 14, -8, 9, 3, -8, 9, -2, -6, 4, -10, 0, 3, 9, -12, 15, 0, -18, 15, -8, 0, 4, -4, 8, -18, 1, 4, -8, 7, 4, -5, 1, 0, -2, -4, -8, -6, -1, 5, -5, 8, -3, -6, 11, -6, 5, -1, 10, -4, 2, 1, 0, -12, 12, -10, 3, -4, 8, -10, 12, -8, -3, 11, 2, -4, 13, -9, -7, 0, -5, -3, 1, 9, -13, 6, 0, -2, 12, -2, 0, 2, 2, -10, 4, 9, -6, 0, 3, -1, -9, 6, -1, 4, -3, -2, 7, -13, 6, 0, 0, -2, 4, 1, -7, 6, -3, 3, 7, -9, 0, 4, -13, 14, -1, -7, 9, -7, 10, 5, -5, 6, -5, -9, 17, -6, 0, 0, -2, -6, 0, 5, -8, 5, -6, 6, -1, 6, -5, -1, 0, -7, -7, 7, -9, 7, 6, -1, 12, -6, -4, 5, -7, -12, 23, -18, -1, 12, -10, 4, 5, 10, -8, -1, 2, -8, 11, 2, 1, -4, -4, 0, -4, -2, 15, -7, 0, 7, 3, -9, 3, 0, 0, -10, 14, -8, 2, 0, 1, -1, -8, 12, -18, 6, -4, 4, 7, 4, 3, 5, -10, 0, 3, 1, -4, 3, -10, 6, -5, 7, -1, 3, -3, -7, 17, -7, 2, 5, -12, -2, -5, 0, 0, -3, 15, -8, -1, 8, 0, -3, 3, 1, 5, -4, 2, -4, 3, -15, 8, 1, -8, 5, -5, 17, -20, 9, -3, -13, 6, 4, 2, 0, 6, 1, -1, -2, 3, -5, 1, 9, 1, 9, -2, 0, -9, 4, -5, -8, 14, -5, -5, 5, 1, -6, 9, -2, -5, 5, -12, 6, 4, -2, 0, -2, -5, -2, 0, -1, 12, -1, -4, 13, -7, 0, -2, 5, 1, -1, 10, -12, -7, 2, -6, 1, 4, 2, -18, 12, -4, 0, 1, -1, -4, 2, 2, 1, 9, 0, 0, 4, -8, 5, -3, 10, -6, 8, -10, 4, -3, 7, -5, 10, -3, 1, -3, 1, 7, -23, 8, 0, -6, 3, 13, -5, -6, -6, 1, 1, 4, 0, 7, -7, -3, 12, -11, 5, 2, -7, 7, -5, 0, -9, 8, -11, 17, -5, -1, -5, 1, -10, 2, 15, -10, 7, 0, -8, -10, 11, -10, 6, 3, -11, 10, -4, 7, -4, 4, 0, -14, 12, 3, -15, 12, 1, -10, 14, 0, -8, 8, -4, -2, 4, -9, 6, 0, -8, 4, 0, -4, 3, -9, 19, -17, 5, 11, -20, 17, -10, -7, 6, -10, 1, 14, 4, 3, 14, -17, 4, 3, -14, 0, 7, -11, -3, 18, -13, 4, 0, -7, 5, -2, 3, 0, 11, -18, 10, -5, -2, -4, 4, 0, -8, 5, 4, -7, 6, -6, 1, 0, -12, 12, -3, 7, 0, 8, -2, -7, 7, -11, 1, -4, 4, -4, 1, 11, -8, 0, 5, -8, 6, -8, 7, 0, 0, 1, 0, 7, -17, 18, -7, -3, 5, -6, 12, -3, 3, -3, -5, -3, 0, 0, 14, -20, 10, 0, -9, 4, 1, 2, -2, 15, -13, 3, 7, -20, 3, 9, -8, 5, 9, -11, 9, -10, 0, 17, -15, 13, -2, -12, 8, -7, -6, 11, -4, -7, 5, -4, -1, 0, 2, 6, 4, -1, 8, -12, 5, -10, 13, -3, 2, -5, -1, 2, 0, 7, 0, -6, -2, 7, -19, 12, -5, -3, -4, 14, -7, 2, 11, -8, 0, -2, 0, -10, 12, -6, 1, 11, -13, 10, -8, -5, -5, 0, 6, 4, -5, 2, -4, 0, 4, -7, 18, -15, 1, 4, -11, 11, 1, 5, 11, -10, 0, 0, -10, -2, 15, -12, 4, 12, -22, 6, 0, 2, 7, 6, -3, -2, -9, 2, 0, -8, 14, -4, -3, 3, -4, -2, -9, 10, -2, 3, 9, 7, -7, 1, -1, -2, -9, 13, -8, -4, 6, -7, 5, 5, 1, 5, -3, 0, 1, 1, -1, 9, -21, 12, -9, 2, 10, -3, 4, -4, -9, 6, -8, 9, 3, -11, 9, -12, 8, 5, -4, 7, 0, 1, -3, 0, -2, -5, 12, -5, 7, 5, -10, 9, -18, 14, -11, 9, 7, -1, 5, -10, 0, 5, -1, -1, -1, 2, -10, -7, 11, -8, 9, 10, -5, 8, -6, -17, 18, -14, -2, 15, -12, 5, 3, -1, -1, 4, 1, -2, 6, -18, 5, -5, -8, 18, -8, -1, 5, -8, 2, 2, 11, -2, 3, -6, 0, -3, -3, 14, -14, 6, 0, -7, 8, -12, 14, -1, -5, 11, -5, -2, -2, -1, -7, 11, -4, 8, -1, -4, -9, 0, 0, -2, 8, 2, -9, 12, -3, -7, 0, 0, -7, 1, 10, -5, 2, 2, 1, -1, 5, 6, -12, 7, 0, -1, 5, -8, 11, -10, 1, 5, 2, -9, 24, -26, 15, -2, -17, 12, -8, 2, -4, 14, -11, 4, 1, -2, 0, 3, 13, -9, 1, 8, -17, 10, 4, -7, 9, -4, 0, 11, -10, 7, -5, -2, 5, -1, -1, 7, -17, 10, -8, 15, -2, 4, -3, -3, -4, -5, 12, 0, -3, 6, -1, -1, 1, 0, -3, -2, 0, 8, 3, 2, 3, -8, 5, -7, -1, 15, -4, -1, 11, -5, -17, 24, -11, -5, 11, -13, -6, 11, -3, 0, 3, 3, -6, 6, 1, 3, -2, -5, 10, -10, 12, 0, 3, 0, -3, 2, -12, 0, 4, -11, 2, 8, -1, -9, 5, -6, -4, 11, -5, 10, 4, -22, 23, -14, -2, 15, -3, -6, 8, -11, 1, 4, 9, 0, 4, -10, -1, -10, 9, 7, -4, 10, -4, -2, 1, 1, -7, 2, -1, -12, 1, 7, -6, 7, 2, -4, 4, -9, 12, -10, -2, 2, -9, -3, 10, 3, -3, 2, 3, -3, -11, 8, 0, 0, -1, 4, 1, -3, 5, -2, 13, -6, 0, -3, 7, -11, 11, 2, -6, 12, -12, -2, -1, 0, -8, 7, 12, -11, 11, -4, -9, 10, -20, 17, -6, -1, 8, -2, 3, -5, 11, -1, -10, 5, 0, -6, 2, -6, 3, -8, 9, 0, 1, 11, -4, 1, 5, -3, -8, -2, -3, 7, -1, 6, -5, -3, -1, 2, 1, 4, 0, -13, 12, -10, 5, 10, -6, 5, -2, -5, -6, 7, -6, 4, -3, 1, -10, -3, 13, -17, 4, -6, 1, 1, 2, 3, 4, -7, 0, 6, -14, 11, -7, 9, -1, 7, -4, 0, -10, -5, 10, -10, 6, 11, -20, 6, 0, -3, 9, 7, -8, 0, 0, -11, 1, -4, 1, 2, 6, 7, -4, 2, -10, 5, -2, 7, 3, 0, 3, 0, -11, 4, 1, -13, 11, 0, -15, 17, -6, 6, 0, 2, -2, -10, -2, 2, -10, 3, 4, -5, 12, -11, 14, 0, -11, 18, -15, -5, 9, -14, 18, 0, -1, 6, -8, -4, 6, -4, -4, 17, -12, 2, 2, 6, -15, 17, -6, -4, 0, 1, -4, -3, -1, -5, 0, 2, 0, 15, -12, 17, -12, 0, 2, -13, 7, -4, 1, 11, -1, 8, -3, -3, -5, -14, 8, -10, 11, 3, -6, 20, -19, 3, 1, -3, 3, 0, 9, -5, -9, 20, -11, -3, 7, -6, 1, 9, -2, 8, 0, -14, 10, -2, -14, 18, -14, -4, 8, 0, 3, 3, 0, -9, -1, 6, -10, 6, -2, -5, 0, -1, 10, -2, 3, 0, 0, -13, 3, 3, -4, 0, 15, -11, 0, 8, -7, -1, 11, -10, 4, -7, 2, 6, -14, 14, -9, -10, 13, -5, 1, 4, 9, -12, 12, -7, -2, 0, -10, 6, -9, 9, 0, -5, 9, -3, -12, 0, 0, -7, 13, -2, 0, 6, -9, 7, 7, -2, 14, -19, 7, -2, -15, 14, -17, 15, -2, -3, 22, -20, 10, 1, -17, 13, -5, 6, -7, -1, 0, -9, -2, 18, 0, -6, 10, 3, -22, 7, 7, -9, 3, 18, -14, 4, 5, -9, 1, 0, -1, -3, 18, -15, 15, -8, -12, 8, -12, 6, -3, 6, 0, 6, -1, 7, -9, 14, -7, 1, -3, 6, -8, 3, 12, -19, 20, -8, 1, 8, -15, 0, -3, 0, 9, -5, 1, 2, -6, -6, 13, -14, 6, 0, -5, 3, 5, 0, -4, 11, -5, 3, 5, -5, 5, -5, -2, 4, -4, -9, 11, -10, 6, 10, -7, 15, -15, 2, -1, -9, 6, 5, -8, 9, -11, 7, 0, 0, 2, 7, -12, 7, 2, 3, 0, 8, -7, 2, -4, -10, 15, -7, 4, 0, 4, -3, -1, 13, -11, 0, 4, -8, -2, 5, -4, -1, 9, -12, 15, -10, -3, 5, -5, -8, 3, -6, 2, 1, 2, 1, -1, 6, -4, 7, -2, 4, 0, 0, 3, -8, -4, 2, -17, 11, -9, 6, 1, -2, 5, 2, 6, 3, -1, 8, 2, -5, 11, -6, -9, -1, 0, -5, 13, -3, -4, -2, -3, -6, 9, 0, -2, 7, -13, 5, -1, 0, 3, -5, 12, -12, 19, -8, 0, -2, -2, -13, 5, -3, -3, 13, 0, 4, 3, -2, -8, 1, 0, 3, 0, -2, 12, -11, 3, 3, 5, -8, 11, -7, 2, -10, 7, 4, -6, 6, -10, -3, -5, 1, -1, 7, -6, 7, -10, 8, -6, 7, -7, 17, -10, -3, 11, -3, 2, 9, 1, -1, -10, -3, -3, -10, 12, -3, 8, 0, -3, 1, 1, -6, -2, 4, -5, -4, 9, -10, 0, 6, 0, -5, 12, -11, -3, 11, 0, -2, 10, -12, 7, -6, 7, 6, -12, 6, -4, -3, 8, -1, -6, 13, -12, 8, 7, -13, 5, -1, 0, -1, 5, -4, 1, -2, 15, -11, 13, -5, -11, 6, -3, -6, 4, 3, -5, 2, 17, -8, 3, -3, 3, -12, 8, -2, -14, 7, -2, 9, -4, 4, 0, -14, 8, 1, 2, 2, 6, 0, 0, -3, -1, 1, 0, 0, 0, 0, -6, 0, 1, 11, -4, 4, -5, -5, -7, 6, -6, 12, -11, 6, 4, -2, 0, 4, 0, -7, 4, -1, 1, -5, 8, -7, 1, 9, 2, -3, 1, -5, -5, 4, 0, 0, 0, 0, -1, 10, 6, -7, 10, -6, -1, 0, -2, 0, -2, 7, -2, 5, 14, -20, 10, -2, -2, 2, 1, -3, 0, -12, 17, -7, -2, 13, -13, 8, 1, -3, 12, -10, 3, 0, -6, 10, -10, 9, -8, -6, 14, -17, 9, 2, 0, -8, 7, -8, -2, 4, -2, 6, -4, -3, 4, -6, 0, -5, 12, -6, 0, 2, 1, -8, 6, 7, -6, -4, 4, -5, 2, 7, 3, -3, 1, -6, 0, 4, -8, -1, -3, -5, -2, 9, -4, 6, -3, 10, -6, 4, -3, -1, -6, 1, 4, -4, -1, 12, -14, 4, 0, 5, -11, 4, 4, -11, 4, 5, 0, 0, 0, -4, 10, 0, 4, 10, -7, -6, -3, -8, 11, -1, 3, 3, -6, 0, -1, -1, 8, -2, -7, 0, -10, 4, 5, 1, 2, 1, -7, -1, 3, -4, 8, -1, 1, -1, -7, 9, 0, 2, 12, -11, -4, -2, -15, 9, -2, 12, -5, 9, 5, -17, 13, -2, -13, 7, -11, 2, -3, 9, 0, -1, 8, -11, 7, 5, 0, 0, 6, -8, -2, 0, -3, 4, -7, 17, -7, 0, 8, -11, -2, 13, -6, 7, 0, -9, -6, 0, 0, 0, 6, 4, -10, 10, -1, -3, 0, 3, -14, 13, -7, -4, 17, -8, 0, 1, 3, -2, 8, 4, -8, 0, -10, -7, 9, -8, 2, 12, 0, 0, 11, -1, -8, 1, -5, 4, -6, 5, 10, -10, 8, -7, 4, -13, 10, -2, 0, 0, 4, -3, 2, 8, -10, 10, -13, 9, 1, 0, 3, 7, -9, 12, -15, 7, -1, -17, 8, -5, 2, -2, 2, 15, -8, 5, 1, -7, 5, -5, 0, 0, 0, -1, -3, 6, 0, -1, 3, -3, -2, -9, 0, 1, -10, 18, -4, -3, 15, 0, -10, 8, 0, -9, 3, -1, -3, 4, 6, -2, 7, -13, 12, -5, 3, -2, 0, 0, -10, 9, -6, 5, -6, 3, -1, 3, -10, 14, -14, 0, 4, -11, 7, 7, -13, 10, -10, -3, 7, -13, 8, -1, -6, 9, -2, 7, 0, -6, 13, -7, -4, 8, -1, -6, 12, -13, 3, -3, -2, 0, 0, 8, 0, -5, 3, -5, -2, 0, 10, 1, 3, -4, -3, 3, -4, -4, 6, -3, -13, 15, -2, -1, 4, -3, 3, -10, 7, 7, -13, 12, -10, 0, -1, -7, 11, -7, -6, 15, -17, 13, 11, -15, 15, 0, -18, 8, 2, -7, 4, 9, -12, 9, -7, 5, -5, 1, 0, -8, 5, -7, 11, -23, 18, -2, -3, 0, 4, -6, 0, 8, 0, -8, -1, 2, -1, -3, 6, 0, 0, 5, 0, 2, -3, -15, 17, -13, 2, 0, 3, -1, 0, 10, -15, 12, -10, 10, -1, 4, 0, -7, -8, 9, -12, 0, 18, -11, 6, 0, 4, -12, 11, -10, 0, 11, -12, 11, -8, 1, 1, -13, 15, 1, -9, 7, -2, -6, 11, -6, 13, -19, 5, 2, -3, -2, 10, 0, -8, 17, -17, -1, -2, -10, 19, -14, 8, 7, -9, 3, -7, 3, -10, 1, 5, -2, 5, 4, 0, 9, -15, 10, -10, 0, 14, -13, 10, -1, -15, 7, -1, -8, 10, 4, -15, 4, 0, -6, 4, 0, 8, -6, 5, 9, -10, 7, -14, 17, -8, -1, 6, -9, 5, 2, 2, 6, -7, -8, 7, -4, 9, 0, -1, 12, -22, 10, 0, -17, 22, -18, 7, 6, -19, 23, -5, -2, 9, -3, -9, 5, -8, -10, 12, -7, 6, 4, -5, 14, -17, 10, -3, -12, 5, -6, 7, -1, 1, 5, -13, 12, 1, -6, 9, 0, 0, 5, 0, 0, -3, -3, 0, 0, 1, -5, -6, 1, -3, -5, 0, 4, -7, -1, 7, -12, 9, -6, 9, 0, 3, -4, 1, 1, 4, 7, -1, 2, -10, 0, 0, 7, 3, -9, 2, -6, -5, 11, -8, 11, -3, 0, 20, -9, 4, -4, 3, -9, 5, -3, -1, 0, -6, 4, -8, 13, -7, 4, 13, -19, 7, 5, -8, 5, 0, -7, -3, 4, -8, 6, 0, 2, 1, 8, -14, 0, -6, -6, 4, 0, 9, 3, 6, 1, 0, -8, -2, -3, -4, -1, 6, 3, 1, 0, 3, -1, 0, -4, 4, -1, -2, 0, 8, -12, 6, -2, 1, 11, -5, 9, -5, 4, -18, 10, -3, 5, 1, 2, -3, 3, -3, 6, 2, -10, 3, 1, -13, 5, -2, -6, 4, -8, 8, -1, -2, 2, 12, -1, 0, 2, 4, -13, 0, 12, -20, 20, -4, -2, 11, -15, 0, 5, -10, 1, 17, -13, 3, 11, -9, 3, -5, 4, 2, -11, 9, -7, 1, 4, 0, 9, -19, 14, -7, -1, 8, 2, -4, 0, 8, -5, -9, 6, 0, -5, 3, 6, -9, -5, 5, -3, 2, 8, -6, 5, -7, -5, 4, -1, 7, 4, 0, -7, 6, -17, 12, 0, 2, 12, -8, 3, 5, -14, 18, -10, -7, 9, -10, -4, 6, 0, 4, -2, 7, -5, -2, 0, 3, -5, 7, 0, -9, 13, -4, -5, 2, -7, 4, -11, 6, 5, 0, -10, 15, -10, -9, 14, -5, 1, 3, 3, -15, 20, -17, 7, 9, -13, 15, -10, 3, -13, 8, -17, 4, 8, 3, 1, 9, -8, -5, 0, -5, 5, -3, 11, -11, 12, -6, -2, 0, -3, -3, 6, -2, 8, 12, -8, 15, -12, 4, -6, -10, 8, -3, 4, -1, 6, -5, 6, -8, 11, -5, -14, 11, -9, 2, 4, 0, 8, 0, -5, 4, -2, -17, 7, 0, 0, 4, 6, -5, 8, -12, 6, -4, 0, -3, 1, -7, 3, -4, 13, 0, -5, 9, -10, 7, 1, 0, 8, 2, -1, 12, -11, 0, -4, -10, 8, -7, 17, -19, 7, -2, -14, 14, 2, 3, -2, 0, 5, -11, 2, 9, -8, 2, -3, 8, -5, 5, -2, 0, -4, -3, 8, 0, 0, 7, -12, 15, -9, -2, 3, -7, -9, 12, -4, 2, 7, -4, 0, 5, -14, 4, 6, -7, 6, 2, -8, 5, -4, 4, 4, -4, 8, -7, 19, -20, 8, 5, -13, 5, 11, -22, 12, -1, -10, 15, 2, -11, 17, -10, 2, -4, -7, 12, -3, -3, 13, -9, -12, 8, 0, 5, 6, -4, 1, 1, -6, 6, 2, -9, -3, 13, -21, 13, 2, -6, -2, 7, -10, -1, 13, -18, 17, -7, -2, 7, -9, 4, -5, 0, 0, -5, 20, -22, 7, -5, -1, -1, 3, 14, -15, 1, 12, -6, -5, 12, 2, -8, 2, 5, -1, -2, -3, 2, -1, -8, 17, -12, -3, 5, -12, 5, 11, -3, 0, 2, -5, 6, -12, 12, 0, -12, 5, 0, -3, 1, 0, 2, -7, 4, 1, 0, -7, 17, -18, 1, 10, -17, 6, 8, -4, 7, -5, 3, -5, -4, 9, -20, 11, -12, 1, 10, -10, 5, 1, 1, 5, 2, 6, -12, 1, 9, -7, 1, 4, -4, -7, 10, -1, -2, 21, -15, 7, -8, -4, -3, 5, -2, 12, -7, 1, 4, -14, 9, -1, -6, 3, 9, -8, 9, 1, -10, -3, 4, 1, 3, 1, 4, -9, -9, 18, -8, 0, 8, -6, -4, 0, 0, -12, 18, -6, 1, 6, 0, -7, 4, 13, -17, 15, -9, -11, 13, -3, 4, 10, -11, -4, 4, -9, 3, -3, -5, 5, -6, -1, 13, -11, 5, 5, -15, 7, -8, -2, 11, -1, -1, 4, -13, 11, -8, 11, -7, 7, -3, -9, 17, -13, 1, 6, -15, 15, -6, 6, -2, -1, 8, -1, 0, 13, -2, -12, 5, -5, -1, 6, -7, 3, -6, 2, 7, -11, 7, 2, -6, 2, 5, 0, -12, -2, 7, -15, 4, 11, 3, 0, 10, -7, -7, 12, -15, 10, -6, 7, -6, 6, -3, -9, 7, -4, 10, -7, 6, 0, -20, 10, -5, -2, 2, 7, -7, 9, 0, -4, 2, -3, 4, -8, 9, -13, 0, 0, -5, 9, 3, -11, 10, -7, 5, -4, 8, 1, -6, 10, 0, -13, 17, -9, -4, 9, -4, -7, 15, -19, 17, -11, -3, 9, -2, -3, 4, 2, 3, -3, 2, 1, -1, -2, 2, 0, -2, -10, 5, -4, 2, -3, 6, 5, 8, -6, 8, 0, -10, 5, 13, -9, 0, -3, 0, -5, 1, 1, 8, -15, 13, -7, -7, 9);

    signal memory_control : std_logic := '0';      -- A signal to decide when the memory is accessed
                                                   -- by the testbench or by the project

    constant SCENARIO_ADDRESS : integer := 1234;    -- This value may arbitrarily change

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);

                o_done : out std_logic;

                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,

                o_done => tb_done,

                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;

    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.

        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;

    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_rst <= '1';

        -- Wait some time for the component to reset...
        wait for 50 ns;

        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench

        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock


        for i in 0 to 16 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_config(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);
        end loop;

        for i in 0 to SCENARIO_LENGTH-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+17+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);
        end loop;

        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component

        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));

        tb_start <= '1';

        while tb_done /= '1' loop
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;

        tb_start <= '0';

        wait;

    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;

        wait until rising_edge(tb_start);

        while tb_done /= '1' loop
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH-1 loop
            assert RAM(SCENARIO_ADDRESS+17+SCENARIO_LENGTH+i) = std_logic_vector(to_unsigned(scenario_output(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(17+SCENARIO_LENGTH+i) & " expected= " & integer'image(scenario_output(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(SCENARIO_ADDRESS+17+SCENARIO_LENGTH+i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done == 0 before start goes to zero" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;

